PK   ��U܌W�Sq  �    cirkitFile.json�[�$9�&�Wg^��_�mgw����b�*ᰛW&:N�](�_�����I2ќ������2�˩�)�")����[�o��s��6��m|������O\z�s�6��~�+�����������_����_�7��el�������J��.�QV��ukdǌU���Sgvf/?���O�S�h
�����Y�1`)��Dc�R`g�ƀ����K���;[4,vvhX
�������+J4���@U�u%�+K4���.�$
��D�(�*M"��+M4���6�$
��D�(�M"�Vx݉&P�u'�D@A`h�u���N4���;�$
��D�(�M"���N4���;�$
��LH�����ּ�������/�_ڷ��	_��݉����������y�V3��f4�o�}��kڞiz/;�����O$���x�4��F��k��l��N5L�ΏJ��3�CR�	�D�����q�mF�F�V6��;����p���		VN@<��8x;�hy�V_Lӛ�kՅ����H�<!�Il�j����1^�^K�(w雠�l�Tk�(���-'���$<!#W�aa�wA����(���S�o.B������Ŗ�?����p|"E�StYy��i9�F�V7J��q��F�ӽ����-�-�I�qZt�iy�iyG��ӢcgC�;C�;Rt�;[Z�YZޑ�����������E�Ξ�w��w��8-�x'C�<��sH��'�o�����9��K����`��K<��%vlh��<b�;(��81�x�H�?bO�'�oM��G�m������}/1��=Z|�_��&���A���w���#�<h�qb|1;����->N�/�5��O���81���A�?b��'�sI��G������b1���Z|�_��!���A��㋙G��#�?h�qb|1g����->N�/f{�����ǉ��<5b��)�l*�`��v��|�Žo\�X�;ێ���0d�������3`��A�����|w櫮w�k�8%t�gM�\���]o��~~���i}�D���/c��꛶m�J_��ڿ �権]aj��}�/�(�J�.�u���7�K16<��2�+���眵^�ˈ%S@�'J�05(�h��a���v~��d��(��I�6 f�!�����.n�,	Ç$�D�!�P����2K��ϸ�A
��L���RP�~������ ,>= CRf)0���@�BR�`��x�R^\�k�����Y
�z���%!�CY���}���G�=�������kn/�_�ȇ�z�y�����ј�t��!�>;���d���V��jj��Zb�6%�4�BM�Zk����55j�-jj��ڡ�昩=jj�R)(uV�~��F�b�67J�)��s�F+�	`s�TZ1N ���N�PJM��7Gi5��j��$N�QzM���^���[���D�o��k��J�I�>(�&Q�E���B����J�	�^SE�6ڱ�ؾ�i�4o�V�f�t�������ػ�E�C��p�!_GmPQT����6;���b���!S�����:j���R�L�.����[����B/{�I9�
�>��4�F�
�}�I�N?��)�349r�&���~u&���	�{]�i��Q�2�5�F�����Zt4@s#�+�p�H��ro{���>�B�ܭ8��kROm��Q���%r�J�n��U"���mW�	�ܭ�[9΢���*�ƬDY��AH�9�P'�9
�s*���q�K����w�0�c��o�X�ӻ�ҍ���u�*�%�8����i�(E�J�2h�P&���\�D!���)	ԩ�KG:h�PN�Ʃ\8N#�Z�$.�U�@k�cN��o�@��	P�ri��֩���'?�F�k��6���F&.>�S�vl������`S�4u�M]�1AS��'l��K��L]��M]ڝ��K�?h�����x���t�æFm��3����98��u�D�͍�g����8 ������/�~�}��þ�<E7�հe�yVb��_��a�G�_�.d�������}��%m1�~��K(lj��Gi\�����Q�eJI��Zr�aS��W�[l��Z���F���k`��(���͍2`��-ln�J+�����4�+F�a�3j�)�VS�=V�Ô9J֊�u�ܨ=����Fp�}�颐��B���fXdi:k�鬑��F��}��i�����2��K��Lf���,v���t�K�`BqȽf�{� ��A�5��k���@'��m��	��DU)^�l`̯��_]�+��5bj�]�E1��-A�z�Ԩ�8�bx�0��S�.�������T�(ԯF��-9���qP�V�Ƈ��0s�4,�WB wp�T���0�N+�"Bo�1g'jj\����{�(9/�<�FI1s��ln�Ը�((�a��
�}\4Gm��Yhd37J7�TS�fe�,��i�^��_P�xk���̍�/(Ն{eaQ*�xm\o�F)ޛAo�0s�tJ5��`�R�ȇ!��i��f�q��7�R-�k3�z�T*�=J�q��s�����(բP6�E�T�[�b��ި����47N���A�R��w0�\u�:f�Q�ƽ(4�.B�&�C���Ň0@�A��e.43w9����r���`�
���O�S��_�!�.�>Ї����/q��x�S���F�u��}���a��p_/�`/���3�`z��r���e��!�n��%��H��xa�|��i���#�#M�}��o�	�TR�7�a�G��F� ��XՋJ�/ZW�X��%�z���d�Co�0OPV�E����sL�>�w��؋W�H"&}��,�y�B�1��-
��,�y�.�����=����55J��b+�T9��(��p�2P��p�2P,�g��ڀ����(�Ƌ�vЋ~��(}^L��Bb&Gm4^L���ǡ&ǕAn5�R�H�C��b\&�+&ŀ�Dc&�m�b���2jrT��b�h�]���re�����KZw5y� "�v(j򒆃�DM^�p�j���'�w������0��v�PCm4�i��g�Gm3����e��Ό(������̍R��su���b>�5
fn��F����(��<�QS�J��o�V>���"1sU�W$f�J����]Ti�^����*�+3wQ�{Eb�.�4`�H��E������Հ�"1w�E�����׊e�`s��.�P�!����@�o\��X���37j���b�hOsL�j�RP�uz��Fmn���(�fP6.�e��v�Ai4�Bs������S�Ԩ�Fi3�̀t��=t�׌KRq�(h��M���_���׷���z'׽��н�o�Y��i%�q��F�U㺎5�cƪ�Z٩�����?�韗O��T��.�4��M��i��m� ""4��ADDh��M�����,����8""BS[rDD��n�4���ЉT$�֦S�dz��)n*Jsw"Ld���)o*Js�w"Ld���)p*Js[z"Ld:��)q*JSj&2=.��8����
��Mg���qA�ǩ(����dz���r�0��qA�ǩ(�)���dz�D���Ʒ���C9����}������o��?�)կ�f�V��C��C��3���C�zV~ְ��8��)V���`egy ��7�x��g�����:��G`�`eg}_�!|=+?+;�C�j��X�!X���W{_���������C�zV~Vv������#��C����C�s^�Z~�x�sos��@ˏA�mΛ!`�1��!h��1�=��:-?m�<���x`���Ǡ������/�����������6�;��c��C��c����cx{�GvZ~ژpo���AˏA��8�/;-?m��8����e���Ǡ��%��������1O������6����c��C��c�Ƽ�cx{�_vZ~ژuo���AˏA�Ȏ��1~�!h�1hc>�1�=�/ˠ�HIʢ%�I:�/��e���0��'����Z7N��d���S�mx�����h}�م��\T�\�˥���\뇶�M�;�(�}�Z���v���s{l����Tx^�wR)d�ߩ��8/�����L��@��9g���2ο�Z5��L�ȶ�:���bZ�ѽk�\�8�|�u��^�^���`'�B��N*UȚ��Jw}`o�u�j��C�]�7!F��륭K�J�/�/b�4��.�KߴCg�ZkG!.�5�P�� Qݍ����f�nh�he�G�4�`���n�D���!T��h��3��h:wc�tC�B� ���D���@T��HA�ّ7\�p�x�V_Lӛ�kՅ���� �R� *�����T74�u]�g�w�a�u>lU!|;�"4��/Q��:�������$��$�SXTe�ZsT&�1��_4�g
f��8�����C�ez3��)Yd��H����(,�~���hzI�Z�t��M����Q�;I�7���U|�j%��$���Av2jFÄ0d&	֗vP��^�/GGC��|huъs-:�:c0Zo�bv�<F��׳�VPzo~����)�ߨ������4�*��\^�Z��o:��T����r�Kr+K\�Ġ"�U[V����A��I��� *�E��TO���ܝT\�x�P)���+uU�	Z�vV���r`���lHT3�@dh$�Txd/[5G@d
�����U���h�x>�7m,)�O�M�D�Pb/�����1dh�x>�7}K)������($�K^��Adh�X^m�6Ɛ��b���)�4����شN�֔4���@dh�a��a�Nc�LR샿+[U��Adh,
5�|`=�hSW)֗ A2�R ���b}��<�2W]<j��D5N"C���kD�K�J׳��o1��6���LU�ַL��	�26*^
��h�x-�
�_^�k�BH *��J5��R���T�G *���J5x�R���\cfT�= �2���ì�5�+i�9�?_��j��Tu�L�������02U�F�F��c02Փ���^�L�������R�ɽdh��T�q/).UM�KƑtKmB�I���G�@�uK, y�ͱ �i7����@ws, }�]c�0���902�����>Vs�adx�ထ5�FF��f]\�����bE���EQ����B�X�Ƣ��`dh�X�H��
����ZF���#�k�1��K#ņF��)64Rl�R�V� Q�5sDE���ATd�&Q�&ҁ�TcH *�vS�bk�9����̂��������j F��	
##j�02U�FF�º02�o�U�Ș��,���9c02������3ô�ݨ���	##hT���7�ad�g%�̢���02U�Fƒ�Psi+�F���N]VsTadx-2##H�9����#�j� ]���T��`d���l:W���TcH0���&si+�FF�"Z02�|Eb��1��l:C���D���0Q׷%�l:���H�CB��z	FF��7si+j#S�'���fE��T#�02�ľ�����^��~l��mN�@����t#���z+cB���"j�D���A�����!T��5���Q���@T���J5��R�� Q��j����JuOä�Hxi����#C#���ؖ��M��F�f?�oadhvT��F�fO�oadh�n�������!���E�a���Sad\-�#�k!:�!�ja(^��ȈZTF��FF�|]]sad��02�vM#�j7l02�v93�X�^F���`dD�h&����N�a�N5�	H�P�ѵ���!��8��nҩ&������i�.h	.hN	^5�CsNpAsPpAsRpQ�mҹ�姌@:��&��w�����t�ѩ�s2M���HKsXT��x��t�`�}y��43f��6zD5�	FF��������#cI|�Y�}5Q��EH�e�`d8��o��jty��ԢR�(��v}+�Ff>:7�`d����%��;#��;#X����F���F���FF����&�Du����#Q��M >��h^�D����hg�Ts�`d�+3g��=cH'I�W�뇑�$^����p�D߸j�������&:������}|��w�����k�6@{r�M�u�������^B���\5���'	""Bs5ODD��ʠ$���UFI�+�� ""4W?%ADDh��J����\���k�WI����6���d���ҵ�-&2��ɔ7�k�]Ld���)p*J��4��t8'S�T��e�i0��qA�ǩ(]&�`����p2=.��8�k]hLdz\��q*J׊�4���� ��T����i0��qA��K���5e����T���T�!X�!XÙ}_�!|=+?k�C��U��#��C���<����������!|U��������>��G`�`egs_�!|=+?+;�C�j��X�!X���Ww_���������C�zV~�x�q�cp��uZ~�x�so�r����1�?��:-?m�W;���x_���Ǡ�����������������6����c<�C��c��{�cx{�7vZ~�x~o���AˏA� ���1^�!h�1hc>�1��e���Ǡ�y��������1���t#vЕ�1~�8�/��e���Ǡ��>��������1o������6�_��c��C��c��<�cx{�_vZ~ژwo���AˏA�����1~�!h9����z��֍SB7�q�tʵoy�����2wR)�rߩ\뇶�M�;�(�}�Z���v�-�S|l��
�B&�����R�����]��.�s�z�.c���T���i9�F�6��r}���]�{%{��*,U2��TF��>���A5J�!Ȯ#�a������R��E�/M�����7��ن���QǇ`� Th�T���q�mF�F�V�}$L3v-o�� ��4�J��j�rM��n�n�]��\Hd��}���T�J��!h4;�N�}��iz�u����1��Q��"��/b��NuC�Y�5jp��}��]��V·�_�R�E *4������A��oz��9�s8BD3����ۋ�A|P�@� ��3�Rx���J���N*�W>;����RxI�Wꈄ�FzKO���������dh$��|y/.=�K�F�KOq��!��4R\z�����^��%C#ť��Ȍv�/�oFf�&�=��Za���u��^��7Q�K�J]h T�2�R���@��B�F^�JB���@RG$�4�8�Adh�pr���H0�����a��"C#ŀ�D�H�H1�����b��"C#�D'w���^24R,i�X�H�$2%h�X�H���bI#ŒF�%�K)V4R�h�X�H�"��i�X�H���bE#ŊF��k)�4R�i�X�H�&r�h�X�H��J�i}�D���/c��pۋ���ҭP�"%�D�*5 *U�Q���JUd@T��Ry�*=��΃I���Ho= #C#��X ���c0242\����Hq= #C��i�������z, F�F�� )��`�.��c02D���c024R\����Hq= #C#��X ���c02D1��c024R\����Hq= �:h�������z, F�ȱ���z, F�F�5�k)64Rlh���H���bC#Ŧ*Ůu���k�Y�x�5�Z�.�S����2�!T��*�� *�UQ�.�
�U�JUπ�T��JU����Hxi��C�����z	F�F��1$�ǐ`dh��C��!��4R\�!���Hq=�#C#�����cH�S�F��1$"S�F��1$)�ǐ`dh��C�����z	F�F��1$"��F��1$)�ǐ`dh��C�y4R\�!���Hq=�#C���Hq=�#C#���L=+jh���k��%}�8�Uӻ�ҍ����� *��(�zJ�JU�A]����!T���!T�/�!Th�R�� *�}�R�� *�]�R�� *�=�:"ᥑ�z�F�F~�ؖ��M�ڃ���OukF�fGխ=�=U��`dh�n����쩺�#Ct*Ј��?C#~�F�,��Y�4�gi��҈�%�Jh���H���bG#ŎF��aBe'QJT�����[@:4;��ﷀth���p�l"��ȶ��K. "y�_s��s��H�H��W]@:D�\���!�g�e'Zu�E'Zs�%'�`D��H��"�C�t�t��!�8D
�H��o�adh��~�#C#���u)�߮���Hq�vF�(�I#���uX��Fn�7�024rS�	�E�h䦞M#C#7�lr�W�&����bG�G�G�G��[A��>��}
��������������/?	����o��/_�~Ο��_߆���?�!7+��B���F��� xhW���W�w~8���?=?3G�,K3�Y�Wɱ�u�6��C�.k�Z���Ni)��*�f`;��g�t�y��U�F2��Ć-$�"�($�� C��:��$�:�vTH�$�*��:�vTH6V��D�xl�B�d�'��7�]���#���Q�D�����	jD�@���#�p�:�r;�V�X��D�!Qd����aF���{�eE�$)a0r��c%��Z`��?lj�PSc���6|�+.5�Y��33��()3��1�Z=A`[=��E��?��{D>��>��|~����E�P�Ņ��CL]^iX�I��*ƕ�S[�K��Z���DL]�p`C���ml[�2N5�8���i��_�Ry�^���.��xޤHPN����ȯ{��@wwݟ�*7���=4,���]�E�0ءe�0׃�_]��07���E���͟�\�3T6R��܆�n�����Y�q���o��������Y�n�vm�L^�ܡ�g1�oX���K�$l�G� ����/���1�#��9^�]Q�/��X1��6<6��35N�;�q���35N���8m�:�q*��|Q�K�f�f���A�a�	0���C��K�0�V�I#a�.�3��E��"��1� ᠩ�wE����O�p��tx��.�к����'��)b���	-����|������|��4��ܺxtB+9"��mo��c��f�i�2�Y�H��:?q�]r�`s��c�7�@����1���)̯.[� u��Zg�VP[75fw!5fs�l]p��ƙ�q������жZ�o청����e���1wQ�B��!�iQԠ����ܢH���L]�D��kPSc'�%sؘ55F���:�F����,/����%�����j�Qmu����$rw�tn�����:>�G7F�aM����+]N ���2T��4�v9�5w)�����]Zo�e-�w�|!�e��P�pw�@A=�n(�������}��r�,�s��>��w��>G����q�,t��>���w���D��1
��F�a��0S���Ͱ�a��U��`sc��D�`bt�DJ��8Q+%@�<���l��ln�f�8Q`��YJs�����1ǧJ��N���{��5Ks��.���_lߌ̴�b�7]+l3\�N��k{a9�nq��˫k1����L-`_:��?p�˪��.��׺��_�d
��D؈�3�9�����;s��6p{"�.�d����?jn��R�A��t�m4��c�lT6 ͍���EZ@s���r�ܨߍ�-�-V��M��j��0����X0�t�|dj�ۋS+���i��^N/�M�Q��QqlǩT�ȑ:��?�s�r�Z-�7�;n�&�m5�j-���{{����T���~p1Lr&����45&���<��tⲧ0	k��19�e���Ƥ��~5&C��M�I,��ASc��O^ASc�˯/a*��K,9��7 �'$(���@=Cw�=��%���O�}��xqn~|�Sc��ӻ��89.;��R֠O�Q�0q�����./ԡ�E�T�>s�'��[�V�lp����jq�Ȅ�������D�nT>*R�P���Vz�sd��ﶸc��l
67�Zf�Yd�%��8�Ia�����ſ6��Kɷ�__�m���!�P�e<�o���.��l2� X�o���=��lA9ț���<�f���<��7����^𥥉e_u{Џ�̉DܠsЏ�ӉDܮs[�@�N< �杛�~DO< �V���~HG����c�TN��jt[�~@��M@?��(q�����G�!�#��FZ��?�B�0c����]���`{��`[�����L_����� ��u��h���츹	���w%��m�ΰ�^�� (J��"�����  ����� � ���v�Ż���� �O.>�m����tm�#�6��# �[>��ϊT��MĂ��o�﫵/�բ�*Qx^č~$�2h���u ��C�-���7�����q�:���jK�5�������1�(,�^�HQ['"�Q�<L�A�-)�>�w4t�� }	�F@}��d��.i��(.`�}��! 6d��n!�>!C�\�
ucm

x�R���6�_����зy���]��h+8E#�
U��F�y ��|A ���|Bs��m�xح.���&���Z��yA�>�g����d#������!5�;�5?�����g��]\����.��C�rӆ�A�`(
0�E��m(|���c�$^9�1��ZOW�G�p4�#��s�<�ZZ��[��l��5��1^0���3a��@ḨR��b 1�J5@HL�Ri�	��I#F/z�	}4�X[�јm���Zm���NG�h@C@h�� }4���4�рF�>*���/��S�з1<|���_b��m��9�{A��hL;���)�BP}Y��`B�HxP:!aj��|%B�C��A��o��ՇM��0էM�� ������� ���R�b��T���(���A�ю���DJ�Ɏ(5e A APJ݁1�A�z�$z	ÃjT��� ��J%� �lG`v#�����JH,���b���t�-/�����=o��7k݃iT�a0}�����N0�3�&���S��>$�P�qc��	�$0�H�J��$����$�F0�"�YLs�j���Z8
��L�p��f���t6ll���C@�*xhS�b���uJ�(h�DL(��11�@d<�6��RM��┬^���c��z)�!T3$`�1�B �:��F�1�T5AC ��,��c$�c)�j�,<�@@��PJ�DP=c���y�C�A�j�M� �IA`�D/�n�	&0G�91g�Y��P�M�@@�f��<�
	Jy�
� I6�F��$��tM0���Q������N[(��̖���( �R��� ��y�c
.������oO0M���Fܓ �( `��j��������Z/����wZ<�D�!�UZ5�!`Z�W�VP��@��I��bZ��g��f��j�5�n�(FC�|���}�Z4$j���8`��F'Uq�l�j�F'I��C�,i�s:Ii,=ǂA �R��F/a�$1ZKKaH�5�9���0�sZ��k��v,���A�jǡ^��~l��m��az�]����X5��v�/�oFf�F1͛��.]��赽���0��V�!�JA� A��,A���"?p�Ͱ�wY4����b-�t8���p�BT����X5ߐ���0�B�/U3�������T-գ�_���P�5�A �������
�Pz�P�������IA0N� QM��B�Q-�$�	�'��`@0��ڭ�1H�F9�۲B��:$Z	u�i4#�6�W��0`N��qkA��QQN��K/V�H4t�$�������4no���R�'��.��0���RB��0�S�@P/h�`�V���1��&ϴ��`�J�o��09��+1��,�݈���V�!�$�W�D�4����e���j�
�b��yP%�H��;V�~���@$u�p��jU>���Z(U b y�Q�'���0����MG�¡�W�ʙ���H�b�����`I�	���$�*ɑ.����:*阆��waD����R�@؆�)u��%9�J��`hJ�c6��酁ٔ��l+=�A QM�4;�?zi߆_?}={o�Ǘ�n��z������_?/?��>Y�6�C�ƞ�8�Vr�w	P�V��:�Ȏ�zke���*맗�G�{Ip<	v�xh�b�M��%�D��E�@�`g�G�&/��(�$���Q�I�4
4	v�xh,�j�B{R�O��	(�Ɣ��A�C9���`�W�� У�@��iL�lx��(S<�)���@�
}��1�[�qPأ)�>�O��<R<}*�)��)�x�T�S<CQx�T�Ӕ�/���o�[��ط?����}������o�{�ǒ��:�)%o0�y��#�C��ܺ�9��{GF>�{�cN�&#�E���F����"���cN��x��qC��}�7�E�|Z|<ŷb���|E�NE�NZ|�;kb�ib�����������'��Ζ�����81>vv��s����ǉ�'�'�->N�/���G���rj��>����À�ɴ95�x�B�����djG�a���!�sB��S#�wX�<��H�rj�������^	1BN�0�R��3!Fȩ�{OjR{'�95�xgK�Cj�!�FyH�#���]91��B��S#����<��S�rj�1G����~
1BN�0�WP��O!Fȩ��jR�)�95�B�Cj?�!�Fsr�yH�#��c>5��b��a̅��!���"\e��x��>�^P{1�ڋ!F�k�O�T�;�n��?gM�\���]l{���nl�$��� r<%Wxy��N6��x����kk|g�1�gˡ+<3�ˠ+�$�K�z����q^����2�l���s�Z/�e���҃j��וJ68����ito�R*�7�:�h�u�W���8Ir�w~?ɽ���/+iAwr��]��tݠ%�$[��E���{is�U��-�\������Z���.}��m�j��p|�l���a)Ub����;K���{ی���;K�f� Z�:��֯}?��/�A��_�J/�����8��Ǎ�7�л��&HEg��_�~�ו^�C�e~]Ao�!�>;�N(�}��iz�u���ޱ�Vc��� r��̯+(Y���T74�u]�g�w�a�u>lj!|��u�ت@n�ׁ���$A��(��b[�%�)�����Kȕ�d���%�J]?`���J���r���:%�i�mRr��6%Wܕ��	9����x�-J�ؠ�oz�}�ӍQ*8mO�h�����(���6�N�Zާ��T�;2��g�n�R�nhWǄ�"sl`�Wd����t�ʋC;!&�P�Z�?JE,�=
zy��(�F�v\�3��Y���
��!l�d��	Ls�������eK�	T�	'�%[�rɋם�OU�-�B����^���-�~�T2�@��<`��d;`��e�	��:����K y���@�m�x�K^_�%�����A
+���� a�:c8̒��H�|��iE��R�v=���K j��C+�2j�9z$V�e*�cGI�P�T��V�X��XkCf��m��7T�v�X�
k<��z6(@�P��V���1+���Jj��$*�a�Z����h�y�����]��q�9zu�<��XR�"o0G�NպA��tx�lhy`��Oa�~%�
؄+!WXM`;��\a7{k%�0�RQ����jE���m�-�r��G��+�+`s��\a[A;E%�P�"��t3��a?�l(Z��F`Ø�ذ�a��s+x#�a���c#�a�`%1��� V�ʌ{	`%1����@j���"���R�6����szd��Ư0z���1�G&<Qj����6~0z��QjZ����cY�Ա��*�И�!��Qj��$��QjO�����t3�Ҙ��E:0�Eaπ��� �P�3@a���h́�Z#k�h�5����J��Jb&�PJ���Kuq)�F/��(OR����������)�<\;̥�CX�>�}�	������X�r���K)���f`��S4A�iN��1=tӸT)]D.�G�
��õо�� c��f���0=���	��FhS҄���l���@��\���7�ۖ�顽����e��ߛ��-�@@��&�ì�V,ڂ<Y ̆Ȥ�0z�(��@��&����>Y �F�E�0�D�J�\�V��`$�����R�������k=h����P(|�H�6���a�7�����<�Ԃ*����˼��(�4��xq� ��Wz(	���yΤ�"�0z��o��R��n��e���f2�J�c��R �Q�ڇ6�N �!Ҍ#^z"��ɹ�l���#���ht��d7��K�5�؏���mc���]w�F��>�UL�ۑb!��1-�8B��SLA���K@��*}C���(}�_}#L
��ƭ������;'��7�.L~�����T,�n�b�6�[ׯ0�}�u�
#��	[ׯ0ؽ�u�
#���-�F ���_a2݂5 S���`��eN{ F/��6sqW0_a�2�u� �^������e�O�z] zw�`���e������%wF/�?P�7B�G�?Jו0�)��ȳK�G��F/s���<s�X��� �hT�^2C�@��2�`�V�Ix枱XeF0�<�Mxz�X�C	f��`6
�T*� �<�F	v涱TH^J H0S �(�g�(��\@��u	f���^&����H0�r)��:����N�\J�^Q�f^y����F/��%3��0z�z�ɨ�R��T�*���e�O`kF�����e*�`�jF	�*O��e�a�GF����e�
a�GF�����e�b�9��Q*	���RH�t��@����TF/S�#��O�"�0z��(��$e`�s��F�sϟ0�+��_&)��=���_��fd�|���a�2E�QA�L�dT�6S4��M��S��?�}`2��1��d
�c��d*�c��˜o���2�f�����{��2Q^�LJ���^�P����O/w:�����9L��姿�@���(���O/�&?�/|z�K�V<�@��<���E�/B��<��Ԓ�H��K��"ɗ �:�/A�Xd��$�~��K<����e�qQ/M��)d<����4�B�S|�4��餟̇iKM�tzMG�tNL�=h�PU�� 5����IMO�uR���\��?����'��L6�dxO��d�Nv�dLN��;<%�NY�S*��pzp7�k���M����F�{��ч�y��w��_�Ɣ?�!Nv��o7e�M�m������wF�7= 30�� �'�L\���)^;Y���Μb�S�p��M!�)�6æ�v�bES�g��L�8��|8�/�ז�m�|�:������-�|w=�6s�Ȝ�1�h̙s>Ĝ�0���=�|;_��*�{�n�����t�4]M�:�U�t}���y��lU}ߣQu����,c��}0
���\5OO�i8d��U���)�vjC�c��*��p�\�s� ��������Y�Q$
��p�s8$�D�s� �1�J��d�s��(p��JJ����q�նk�u���d��[:]�Q�jg�,`��T��ʤt��1g�U�O)���ݜhlF�K� �M8�Ϡ)�}`�q��Q��Z�3X)A�K+-�<�ASZ)h������ҹ-Q�<�̞ҥsZ��y4�=�K��<*B�s�SR���8��*ichq����&/�Z�ڮ8��J��+hiX���q��Ky#�� ���e�F�lt��R�
�tE
%ʥ�h%�J�K93��
	�:�K)7�2�QZZ,h�dԅn
��X��Ш��NI�@�^��8�$;жިt�N��v-Ge+�pJ� �);*�)�S2�-�Q�R)�r��ؓQ��t��РҖDM9�@�J���*�FF����BF%�e/��Ǩt��:�(u�J��ȍ�ic���H�2F%�e�F�t1�nΝ�(e�z�,3�O��1*�X�g����s��Ҁ����)Q*��)3:P�t F	ʜ��R���r�$�� *=(@�AT:��ؤ
�Q��*��d��UF+����
�e�@��h�����@�[������=�&a2��V��&s|��7l΋J�O�Os`seԓ�N�46�F�8O�Os`ssԃ��-���n����)��F�A������!pP��D���E���z��9�lQ'��jdԠ-*e��%2^�EieT�TdԠEieT���(�����S�8��A�с��Q92*С42�>C���q�r١42��Z.���T2*��sG�C�d�w�sg�C)e���s��Cie�sd�;%J/�ʉ��9�p�Wq+sRx�nF��๳£�s���"Y���K=��R<(�\�*����Ae�a�vx�;��&T�ό.�%�m��|Jp����<Lv^.�	�&�Q�y�D��e/��z�bФ'/浃Р��;�_�РZ4�;�_݀Рn�g'/�a�i?T^{j���UT{�wPڸ��\8�S���Z<9��42�!O��y�*��OF�ߜb�/?36��������RhCQ���)>&��dMg<Q^|	m9��Oj����Bhi�%[��)>-�QD��98(�lݐ�A�fTc���UL)�if�̹U�(��+�̩UL(�A%�Рt2.�=����08���wP[69AF)d\%��./��C;�#6VFsʡ��p2�g1��'s\�ʡݥp2�W1�ڬ'c��ʡ��p2j��X���c>�z�������/�.{�'��o���ӭ>�׏t���~dҏ��#�~���#��'MM9�GS�b�_>��gb�L����3�BY��~�-_K��>�r�L��&��|�ϰy�J�vcJ�ZجR>녢NIꅤNi�_:e�^�S��c:嘾�^��pE�\ы��T��"}:?��E�|Q�bQ�bQ�bQ�b1�:���/4yJ�/4yJ�/����O,�t>���H�]��I��bYw���X�]��.^���b�Hy-���/b�H�"���/r�L�"�Ȕ/r�L�"o
$�\�"3d�L�"��.��.��.��.��.32��v��v��v��/�oW�oW�oW�oW�S(��f�Ϥ�e>��g��L:�Y�3��^����v�2h�u0�:�eLf�/�`�u��:�t�����.|�)_�����.|�)_�����.|�)_�� H�b�ؔ/v�M�����/n�K�����/n�K�����/n�K�����/n�K��n�R���ť|�_|���ŧ|�_|���ŧ|�_|���ŧ|�_|���ŧ|�_|�3!�pv�!�����5�-��fF��7�fY�K>��},��Y�sO�Շ7�%��7{��f��Cw+;5��3;����Nm~7�SK��m��h�w�8����2NMc~7�R+�߭��L�w3)����N⩡�o�O-%.�Hʡ���S[��l%�K�f,��Z�7k�����K<����^���oO-&~��xj2���S���l��o�qm�|9woc;t���p����z����{t���rE�k�����]��j��ȳ8��o������xys�j5J�|�qJ�`�a���_��_�G:����������_�?����/����q��|��������>�S��_���?���o�_�q;Y{�~����������������ti�|Ç�Ʒ�������x��������m^~z��
�k���Kۿ��6�m��q���5���_?����:��~	U������_C��;q-�����F+qR�i�f^������ABK+��:�sM/U�pi��ng�}�������5:���~���v����O���~뿌ׅ����!j���Hu�R����?O_�_����������߾�����X�4�xdHP��v�	�ħF�&8����?2ö�y�~F��%�D�T#������b	3@�b��r��D8Gl����_��'g`ŏ��VŁ.LP��_�����̓�bC��߾��Ňa6g�9�Kdη�M�����>��=���]�%�ve����7���'/4�z��}���׽���m��k�X�q�ez�Ge/|-	�~9 I�fO�㲨ORA�����j?�ON�=5����@I0l��[�=�����i�19�?Z���/�����_����&��$���N
�UA�(L��y�Q��7�Gv8�F���l�1�|Aֆ#ӭ�	��j-L�%NFE�*LT���k%�|`�Q�����-��4nDйF��e8��?Y��6z8{�Azv��Ӹ!��ލm�������K֭��Am-$W��n��7��(��� ��_�[�h�{�ЎS��8yg�3�,��^+x؋R?
oe�������xo�����Z/[9��Z@]� G�p�A=0�)��I&��4��������[|�H��x.ϮG�4PFa��4�X�p_�}��8�HZy=�>E�/Z@.��Moy��� �}`��A�Jvi,��0�1x�*�� �� ,7<�}r:���.�Iś��!���v'�8Ӝ�46̟�Q��^�S�H�ù$n�v�R���`{=�^/:��K�s���w�`���\O�O�GF��nŇ_�L��?.�FYg�c>���|_��=�g���].Ay�6�s1,Xc.^v<���b��5fipâ���a~���ٮ����O��O��n
��h��=�y�g�\ث�$�W�/?�����A7zluPAh���`4��p�,Q8�F� �P]��/;	�d��?y�/�����{p ���(�u1��x��`���<�LpS/���Ps��4ڴ��w�u��]k/�T�E��%\��0X�縂W�����Oo��(t3��b�00���K��)��|��x.��v��r���2P��AM�hoJ�-�J?V؉����O���?��9�i����81ӻYp�qS��	ko`~�����Z�8p�^{�@��T����WM~\�/�a7_��e��*��m�K�ϊNf\V3����̸��ˌ[��=�xV�'�{�������b4�@�lw��d�C��K3�BŸ�i��dp�S�k/d�Q6$���5�HS߭� nj!Լ	�����&�*n��;f��5}��Y��U]8�'�7�3q��e�Dv�LB�ԥ��ȍ��j�i�5�:�u{��[��(3LW`�n��s���K�� 3C�A�iZv�a�*���[�1�q9��q)��0}G4+�`|os73,�g5��<�ܰ+?Auf��@�q9D�q)��"�g�Fn��ܰ��Nv����*��&3,�&7,E��󪟖Q>@�2��S�j�=�
Ы�ܸ��xv����nR��r�r���RD�i�*.)�7!&\f�M����0W`SnX���ۛa)W�r��`eǥ��ӥ��|�k�b??��}���`JG}��1g%l��(�xg#ݛ��A���ŋ�[�5�롹�X�8���j�l�� ��$���.�է`]Nʫ�.cz���_�<��?C��P�&�#^}�D��1����y��WG������n5n\�;��/G�\����~�n�nB�ݢŶ>�̜��q]���������%?"eC~\�����K��Y����+����츌�e���6;��n��/���M��Ӯda�5��\�w�����Y�rv��r�ٕ���r?&;0Ý���3����츏������(���ɏK�a~����Q���L^22
<P��pzԖ��sz67�AE�d�{nX�p�{8Vrr'Rf��Y��<wf���̰�)�'�J#�!>G���Y�|s�.&�.zB:S؄��u�Z" Q/;/ŴY�ŁF���R��Ǖ*�^�XVM��RD?��^ET�#lP|FG�������F�$�-��7v�1��;ܣ)�����ML��ɬ�>d:����0�f��eB��ou3����C��4�
�f�W�ͣO�?Mϙ�ω�\��,�㓿_�������|�(�/�\��
3$/�o�^_�Ǚ�u4�%��'&c�����ӿ��ό��oE~���������g�e��y�H�<Ϟ�9?y:,;�rSD����w�4a���)_��3S�e��r5CaN��v���3��yt��Y�kd7��"���#2sV��� ��4����a��WZ���v��}�=�����q���M��M�dQ�dQ�:��(�Й�M�G��Av������܀N�����)���Sq�����$�6��^5,RX#���s�%�8oT�]�:qi�e��І�Ag�&15H�1X�_�2t̛��D��5��w��s'�nw�֏���w�O<���:�LN�~���i�u,�,ԉ����ֻ������0�Ճ9e�8豑��A :ٸN�`(��Ƶ:�TA����º�oE�7x.z�j�yq+�`0��@
�pƥ	�9i��Z^��ht'/��+��s�Z8�2��8�a������%cgJ�an�CN\9��%f�nIo�[�+m��8�?��?���/��Մ��Bqs��阯��r�'�*P��o�}�x�?VG^Iay�;	ǝ��Ǘ{�%�ݻ>���r�)��>|��i�����ߔ������^�JK����c�c'�rE�����d��t6�aL�뒩�S2�͇��EēE���Yo��)���"����I~����_YLT`��+����x1���a���`⦡&���v��4�� �Q��)�SΘ�%;� �j�2��ǽ,k4fep~��� u'��#�ۅ-�A��˵����}8�|yO��"bsƣ>E�l�����N�q��D�ܬ�xA���W���'��,�Rq��	-��R��q@0#�3S�%���`����	/�&2Ȋ[���$W�&�&l ��m����ό��p���<�}��(�^�ea��j0�l�9�B�t�bA♼m4�M�������I�Yn7 	�L��q�"T�a���"!�ԱE�����N�Ӟ� ��B*c��zc��Z���>��U ��~J�9��I?��O^ٺ-�'�Z��������+.�B��nL�� ���V-�<�@Џ��V��'����U�7��;KH=ɿ�z^����$�o��0�2�x4�J	$N�u���wȆG��Y�q�;$��7�;����f�s��C��T]X$sr2�����n�����?��vN|�t8ab&�Y�L٬�\acF���\��v�7�~�1&d���ʬ Aj�v�0��k�n?7,��	��0�5�,J�X���h$��P��3o?8�^��.H�U��ā�b�?��j|:�.37���0�5�7�E���T@��%f�O��gf&i���Y���,�s@�l�9A*��B�2�D�p��o���6!gw��oؙ���\X[��ܢ�U8}d���S�D�	��k>��sz��:ʍd�.k1��Z��mͯ���an�	+<hŨ����EM�:0cMp�O5F(�e�D���k��v��	�-YH� 6&PK  0K�
��G(<������SP"vV�A�h%آt�l����H��6�x��=)9�o\#���Z̜t�?sZ�`�:����YrQÂMnu8]�KGy_�h"=�q�����%�/����q��d:\����PyX��K�7����I
<�l�����p?�ˤ����Q�R���Y̸�pA�:#ł`�#�J���Ƃ4&o��.����*��v����<�^�Ѯ; ����'9Q������c�M�'!����`p����s�C}�<�����q����$���VUE�<��}$��>��$x��͕�2"��7=XYtg�8�pκ9�$f�_�I�����M�L��).�}τ]�xs���.�wP?��Ӓx|��n7��
���˗��r�D���p���ț�2m�x�r���x��E�3"����X�ٰr2�Uv�(v9��&W�>�����5d��b=l��:�^�ÃEld<w�]�I6�"�Y�EX�������f�p@πGMp׵��87I��c�^�����������b��0k���f�'Q;������*L���͒��?,�*��W�aa���$��s5�k���u�b���i�����*�M������9������c�Y<���8�V��8%��&�n~�������q��xm��q�/�BJ��6����|����Ʃ��_��ҿ~y}���O|����_>����{���ϟ���0}�)�)Br���_��_^ߚ���3����������_���&�o�o�B	5���ǡ������n��<�����ǗX��.�?��)��-���?��?�g�G���7Q��O�a&?��g�ג��=�������?��-�棔��?L�J�8J�~y�F,e�@)[�[	�)e�a�,:?죔����io��̺�������إi!O�I� ������ld����!7�<�-H�{5�ꅭ�#Ќ V�b�f���xR3��B¤Bd�5^=9�達K!��g��P	���G�Ȋ���U+� G�4 VӞ4���;�#O�4k�x0��K���9���"��I]�*�Td��=i����P��~���j,�DW$�t�մ�B<�+v@=F*��JWRq����T�u�R��LzV*v@%���R�V��?��Jb��qQ���gI*�Ye�J(�;�bUu;,$.8t�8���T&�-�t�:"p��
#wo�o����ZS�p��0�1����k +G|*�g8փ����
�hv�l5�$>&e&e�2�@� ����g�;�
>N���|^�t���z�.\�k>��M�#�w�գUgφ~w@=FО=2�/��.�z����+A�+
���	(h֪,h��,gm6$�NRU�.	u�ڃ�(ZO��)J��ϫ'�]���e�+_8�&GqA8Ze� K'�Z8,�p��C���l<2�{#�����F�t� E�.d�ڻ�.;�$c��G���sl��=
x0��
;%���P��>�V�b��tX^B.��K)![~��%p�R�󟃇���^����{��R��dX^BF;KR/DR]��x*";�햐kU.>�c5��8L�c%n�a�x��b�px:����I�C>g{��E�qPiŕ	��O	�5`��|	3=@��Ă!���x{�>V�+J�jTi�%Lg�gt�ӭ�uf%�� ��R����o�h�j-n��jTi���,h؎�7����̰��;��=بD�)euDxR��Y�0�h\.fT�T4���{�<jSCV����ۛ��dQ8V�
��@"����cG�HE(�'������[�M�X�*,����|#px�}M'��{��T4�S��~�h�F]���~Fk����րݩ�Xo�E|���^�r�IY+,�����U��Z�;X��\o�/U���+�ڛ±VXv���q����^�I�$nІD�sэ�"�e�X+� 0G幈h��'ʈ(�K}ʉ},�_�հ��CD���)[J�P�QE��*ڐ�zʁ��bS0V��
|=��\�����"��*jVцD�S콋ȶh<�'>��!c��	�J�
a<TS���6 ��3Co�gئ`<�/�c�2z�����`FC5��h���)��ֿ�o
�jX~�@c<u!�/�G	�n���3���s.������^Dߞ9,�)>}v;��=� ����c����Mب'd˄`��������w�{�Q��~ʄH�}~�)�*�j)J(��z�ZX^w�� ����� ���pd���A������E�?�X�E+|�cQ˭�nU+IWf���Ǘ��j՟�%�U�_ֆ��J���4�y,x�a�׎�T;[aN"l'�H���l�?���^�����2���XM6�^mv{�{w�hh��XX��Ur{5ڃ���ϻx���!40��;=�.�zk�U��� ��b� ���v`�Zs��{�d��7Z��G����3pн��3~��ك�
�T�1uG�g6�5.�~���*%�C�n�[m��6:x*,���[fS�/���î�\�����?�c��X�������3�A|�����Jm���N��î����s�a9�s�>�߿�z(ԟT��9Zu@�3�X4hCwWxX���N�|{�a�Z.�ú���0���[+�A�@�'�)';����S'�h�Ix�76���m�C?�̠���/���E$� � m А ����ʕ��̨{k��Q=X2�Jq�����aBGmk�F	����M�W��Z4@���uEc�SDPR�!j[�6��Hl���p�>~�Z�lԽ���Q=�2�
ʀ�OrtԶm�ё���\�Ԩ{o��Q��[�Q���X��Tm��{��������� ����S����zǨ{W���gW]"�B�$u���F��s���.,��V�����z켹e��\[&�$������۵�/@�+��Ǯ��1�]Y�$h��� l���$�L{�&�3����NI$6� ;����nK�g�ΓZʂ�T��l82	z�V^KP�r&� ذ�t<4m��7u�x[�h�w�����;A���xk���$2V���ްA����z��I�a�ORg�
�H�|.�w-C�K�D�`�
�4}ߔ��A����2���#l��$u~���H����e({��lX���*<4u��̭	V^Y�A5#akIx����pd��\J�J�
wQk	#��b�X�8*8t&�^Ԡ��%a>��N��	�<ʵ��o�A�#4fN�+%W��M�g�-�"�h	[K ���ڠ�"	���A��4��Ihn�㥭�'/�gN��Ǆ�%a�\Q��m�\����n����Q
Z�u�a��'����k�dA�+6�"آ]3���(��&��]#L�K7r���+`6ڱ�ؾ�i�4o�V�f�t��cpj.�{�Zpl 1���h/���֣ؤͬy\s!�<�FԵ1��qu�)�F��ϕJt�@N�W��5$�d)�����%OGT��7�tO�ب����3Ν�����䏃�[���^m.y2�����0��{�M��Ȗ��[S�O<v��[��q����u���%OFԗ��;�����,��ОXU̟��ƠQ"�GP=
�Y��I�Ǌ��j��Sf�j��ucT�Υ�\38ʘ����ʙ��6L�F#����ȖS�C�'v���;�Z�8*(yk��5��١Ӥ�Nx��
�pd���1�^���ݨ`�Y�}��Ώ�'i�sδ.<��,Fc+��/F�r�մ�]���N�X���Q�s�k�X;Қt�v(0��D��lٟ�D[/����z_P!�Vp�a�X�H�FŴ{�0T�^�ރ/� ���Z$��l8*!�5�^	�����BV�O�e4�k�(1�"�k�0�.�� ��e{�$v�#���$VB���b�ߔఒx�9�(���Q�����W��N�I�bOTj82!z���J��\�UpXQ<N�8mY�=sV�m�W�J�o�Ğl���D�l��]�8�],�a�@�Ik%���Bc�hǴ����J��ֈRQ�ˈ,
�pْ�!V���%"m8�4|�w'��Z���J��z�{����F���2.}.�P��p�\���yqb�+^Y�}�T!l%�
�8mtTP�ɸ�7��Ez,�uO�r���
�^�]UTA�G�%����^	�g���[J~,�d݉k�}%'s_	U��N����1�`����k��yؿ1�M9��d�l-Ɠ}{�﫟
a*�SL�X�KL�PV��I��r�Í8q���Y1�vO�Ĕ!p��%q��\�R2{���ݲ�ף̺������/��*b꾍u�7�S��D�+���W�W��
ZLB���#���=��'L�6����F��#|y������%�89�����+h�o[8y����.T��|�)�D�Q%��R��*p��$��Jw_X��Hz�Gʩ��B�k!����BU��'Ÿ�۷-��w'����|�}cA�D*��r�wD��`�Z��qk!�*��S0q��G%l���d��g��j˂�<��<^.i������J�
y+�*��������\���UhA�D�<���6{�?�_Q>Ci-D�Q�W��$��N��po��ƙ�Y`�jA�S�w�p>���.�Hʧ6�E6*+"�5�_[��p�O�8]�?��ق�Ա'��v쟺X�O>!z-�Q���<���-=7 c����W��D�����8������ �R�E6*�\x���Ɓ�p����-���M�n㹫�� �`�E6*/���W���0&�w,䵋�}UlAKD��kWI����"6]x����@���!Z9@�[�ĜT������i}�D���/c��꛶��طB鋔#��ԵN�^w��#k�&�-V+`V����h[�� ҳ�N�QE<��gWs=Jo&��a��w��� ,�c��H�ld��T�p��ߒt�GV���h5(��΂�3]`���;��F&OyNv^'�7ec=����8�SzcW9Y�a�T ���܁�J6�����:	�)�Q�E�0�����*�������#d��l<��u��-x[�dXa�Ls��4Ǯ����]	�ؿ�7�lT��\k .ļ�n[:��
�.`�C<�;v�Z� �ۅ��}�ld���m��R0�FG2�� ݕ'uǎ���%6�ؿ���lT��\�g�g�`�͎dX~�A��d\.fT��)�aqz��Xp�~���1ק��oK�zX~�9�P�O�)��cG��3a̧�c�i�{��7mb;ߎ�ec=,���6�s'
g|?�1�G��|�=ਤC?�n����iE�X˯;,�����3G�9�o�aܧV�7�{�=���^S=Jґ˯�����SE�1��=U���#��{�L��Z�k�?�q�d���=���Qv��@�p!OZy�+I��
��8O���'r��\<�7�����N҆L���Z�dZ�.�ɂ�{����(�����܃�N.�Lf�����N�[��ʷ1:(��<tH,ja�2�R�hW�v�)3���݃�N*��zA:�<jwR�ig��%o�����B2��X���Zʹ]U�a�A���=��������*��bU�B��Nw�՜�ܟx�3;�X�[]yݵ��;��9�{r6�������s�d4�(:�'gҭF-
-��21�T0[�=wU�������؃�N:��h�.�
��8(��B�X=�a�9q����Q&�Rײ�[�cGy�}5�Ǻ��u::�x�Ŝ���AAO��0zudH9��{F� ,��Z�]��a�'�;R�������:]j��x��ɺ�������(%���$l��j�l�%�a9r�ޫ�V��yu�i�v�9��)�s����4�q�g�����T|�]��a�'�a���.�{No8��X57�$������`;�=���k��������<���n�ۑ���d<פ{���<�*����dc1$�c�`n�ZͶl��?�b��OhO���I�!����Ҫ��G�a�$`�D$�6��U�y$��;� �}���X�zTi���IpB�vq��Q�L�UN������;� ��{Zk�>u��p���zTq���
�LE6F������V�\�(��?��e�օuO��N~=�Xi��:t�H;��Ü²V��R���~�N%y�jAi��BU<5.�ʲx�֜�݌t�aE�a�EK5Ԋ�ӆR�s�f��� H�Q�r$Nʸ�����ʝ8S�\k'�
����]�J1���%$�If�ћ����b��V�֋�7����Kx���&�M��)�mld�sɮ����Q�@�L����c����0�E���N�D��Ȧ�d���ǥ�FC#Mƫ��AVZ�?�o]Il1��v���)[��2���p��`�G��y�+�<��3��M�X_������ㆵO� �0��Hpv���`a��k�eG=��� J+���~����sg��#S����ÊM~�b�ZO�&�zL%rje_9.�־�@r`�!�h�^l9�Ê�3,����dE��>�$+���pI��=�E��ʊ�U���B�,I�푾�������8�R_�4��Ã�V25���68�u؅��j���X�cϔ��?���@n v=�9CM�!��zY�sej����k��ܭ�w������ۏ�4V�%_���k����>���}�x���6���PK   �R�Ts�7+5J  dK  /   images/6c71542d-16cb-4630-930f-71c4de5e1144.png4�4\�����G%�F���w� zｷ�e�D	QB�����+��=z������]ks������s�Q�*�xؔ� O^NJ��|��` �_Q3?� y)q���m>�Գ�LWm�5��G8�� ��0P�����h(_׎��hx���๓}��2�Y2���e�`e�e���Kw*�/��|b��G��,�\*k���-/X�F��fg��œr�z�cvvJFK�G/�/i�)m�b]��8�X
�LTjYx�*?>��98����O"2����.d+E]r���q��JW���5,�3E�G\w���_����� �Bĺ9���� !A���7�D�L�2`qx�^2b��z�-|�_�Q��o���O���|�w��o2r|u��؁�P,$,��~��v�7�5==�ʕ�����I���1�B'x��G��'�w��*��#N����G�vW�)�S�J�К�V�%�0�=^뽌�S�13�E�j�^Tj�i�xJ,_3��������T��ٞ�Rd#%*1]{<�+KSH�������`)\�}�^�X&.�.C�f"��#Dj@���a!�B��L ����ecŇ�X�\_@買Ox��-�C�����?����dʲ�J�qQ��s�JC�е9���tx,xXb60u	Ȳ�l�Lˢ�:�l
�Ð��ق��}ǿ��Yn�x�t�E^�M��x��-G���M��άG8�jε�:��C��#�,t�H�M�Q~O���Q�)��%#�!���2�cS�!)�����k�l&m��%�� X�)�t�琰X2�_�N��DE��W�������(�]����R��TI��F���Q��A	�
��)�)/L�<�٣�п��yR6��n)R���D'�-�G\
���FF�K�Ă@g0�/"��9�	�M�#'�9H�a�
B�X
w>KF�"	�|s��/iIġA���a>)5�:뿦���[:y"�B"����N���/$5vq!��}�Y$>��X�3�CF1�y��h9�T#���!� h��+����ގ\WggЙ^�E�-����]�ȂrO�Q�����#���:NSA�Q���|Y�,	�����Rj��[�W����vHpc�z/�4g<QZ�v����&�^�Vɭ���a#���(�|�D�<��MQ�KO�Ѝp�/ �l����Ѝ �d+��ྉG�O��Q��{��ڣ��u6\�@B@����0�g���㒒��QF��c��
MHBQO��3�V3�rP�� ����V��J$���fvf�����v�Y{�{~�Ű?�������E>�=d
�=hh����I���Ě��$�/����š�6�:k��D�0�U;��`�e��gV71"�qq���O�,�ظ������;َۖ�E#�3�=乚����ԭ9LZ?�˾nP�6��e=F@$���'�����`B1@���a��C��4	M(���g�1�Kq��t�-_��,����pV��7$��铂��u��)��eɌ����=���m�������II(8=33�Q~�˼F�~�/�g�K�PxPI��y�6n5[���i���X�O����ߑ'���'�à� �����3V �
��F$j�ö}&=�e(!��s��M���&8���(Rjal#Pi�4���O�>%�|�jm��7o�s۶|�-��w�}�7���aގ9��xh�r-�H�L����=<ʪ
@BD�j�C�r޾�5ȱNw�#[�S>Y�b�I��������V��[���|�b�����=_�kX�Á��FpI�����V-��-y��B����D����^L�4-�G*L����pz�1��
U{�^��6)#g_L��B��['�D�Li:�aAU��ɚ�I�I+@����ދ�4��ޑ�-��؎��M��L|A��"�É������ҧ��T���}*�#O֪�x���ٿZYZ�>�$�������~�<lc�w���]��TW�Z^N0�ZZ2�̇ȧ*�p����;Sc***:����hkk��^��?�%T[��;Ș�������k��g2*Q�����I�ʲ�I�H�(�D��mN����7���X�j����M������(���Qn4t��Q�����}���������@�?�̉������;��&�wڷ�����ɰ�I�m$���2*ʠ�:�Zh=�MX���e&���C��X7 �Kz�G���O#����６|���������m/?��l�"�
tIr���$=�е����_��m���C��^Ӷz6��+^���-G ���%�"O���_鱧%��ώ9��r�!����d�; I���|8˗�(���8���EF��׎W{>��Ńl2#֏{��^szdM�FD'1i��	j�V>�*)Y��yq1��8�	��?I�Qz�C$:��h?�􉅲�_vb/�� b?��m	8*�䍳-������@�{��z���ͪdԹ].��;{���X/V��_�*b8OP�(j������̱K�w܌t�Hjz�:�����Ҧ�5�m9���O��Z=,��X��\�����}�W)m�����CKPe�PS"�N��Jq?WgG�v��kt^E�} ̩����$�R�t_2��QRRv���!tZ[G'x�G���| � ����˥֝�ʳ/5���XP��R�/x(&�ݟ� ��xJͣٴ�[?n�|��ܪ������l�bZ���;o(�5tx�b�x3k��I�Q��U��c	GD'���!F"�Є ������}���8��BP����4f9e[w�o��@�l�&��E�1��p�˷�HQA�ֲP��S��P���n�"%R�Q��\ڐ	(��ۘy��3������Ue;�?�u��)�-p1w�s�Dh~�	���:��;J�VF,FR�}�B�.��Z�Q�g�9���O��!Mr5^Х*V�غq�}�g������d~�xA]����H��ː��w�Nf2 c����R��l����m��]���oyےV�:���i5��D9�1@IYy���X{��>ӹ*����D|��w��¾6}k]�5a߾PI>!�(��B�d�jg��/��P�U��\���l�!v-���1�~�{	C�����7�tp��ফ���T�|P��?�DL���QSS��8bBt嶫������~�������*��[�8]�Ă���$���[m'��4�:i��zP�$E�o�/�2&�������Х�'��:E��,�������l��H���g����=�*������3ܹ`J�`�5'���cD�rN�k`��[L�p��& �S�kV�g��� ]��^Xˠ�;�#��G����4;<��ߗ. ���\ 4W�	����2K�n��vd�L.��x�����e1lC�~	vjЦe'A>s�����%��X������	�+�`������S�8q�Ý~�tgc�܎묎�������[��?����OMu`���3�tߑ��v��۷M����}*�3��Z����K��n��9��d1��>6a����\���YZb�Y�閙�%�2��td*���%��p鈈Q/�����R�_j�HQ��%����k�`�Xo'�VͶ�Gn�;:�+kD�<=�̬�`Lj*���&➞~���lUW� ����4��������*�2����m�������vH��"
��UI!e�N�<"ȇوHq�^��UduW+}/	yo�C.A ��ل(AS�
���+���h���J���}�vCF�!ԓ�H�a�ޤ�;����HRS�уC7���rMC��a@F�,��@urzH��Z/�Ns�gK\ۇ˵�.v����/�4 n�pr&&��DP<�<�
�e���5FO���3UТW��U�~�m��� m`*������z�eˣ�g�>�GF�1	w����o���smJ�M��"�?o�u&T��2&�OؘT~_�=�>s�Lo��K)�<��{ӱk�baB ��TC{���o�B@}�ıi���@�FEa��Q V��ؓ��f`�G'&�LMQ�HOO���`���.�é����F͹�F���F)ju_6��4,P�<!A�e�2���m�Ȼq����4e�����%	MM �� �&�Qr�G:�ذژD�K��@G�ϝ�R�u�+@�#�i��b���Kf�f��M��[����=���q.Ȭ��z�y���9tU�d\ò��pi�xAj��-@�'ڟ'f�	������g#m>���J(�P�:��� '�p�bJ��$�9��v���I�(�����ųv�w�^w�77��1�(��Ǉ�������ՋY#r�J^� �����B*cTlB���
����7n����_�?�;oOM�
|8�ո�������BWM'2�bآ�l�C���+Ε���|�����H ؎������X;ݷx�.L���S.@-V{"L��!���+�ao愯i̹(ҋ����F���!T��z���<�l\U��?�� &	����7s�	�'[[[+�(�N���Kآ(9ݣ5n�|�����ݍ�F�o4nXё�̩�JJ�6�pL�I)����-﹠o���ѿ�ҋР�]w���]�oxx���΅b��w�Q��\`��5^�lu;�m�]��nr�������|g#u5���J�|��*7�\^�4	������ Ȳ��_�)��lO$�=�>��3�q$����������9��ZT�Z������^h�?�pV ��uϝc9f�铀IA�#�� �<J"_��"V�L{Է�o��6"t�A'z�#�}}j�Y4�&���,����Ö�Z�rLB�t�;��r�m��� ��4d�����>i ^d�{�}���H��!]E�Y���]�499���x���g�2�����H� t
y�f ������:��Z��3%"
�L�����>i�>�T����������5������I�����������T�Rl�i� �N���W�0 :�jjL [z�&! �Wt<�ӊ��M8�"m$����g}�@�d��N�?�:�	�2��p�~3�=K!�S4?����giee����wfQ޼u�Vi���l�3�Q^'�X�r��PN���F�ÁE՜�z��@h����v\ta�:��RaȐ�V��Ac���*�'��q�l�d���l����2�*�����}���J����(���dA�镑L�F��-u��	OX����,���ud%#�x
��s+b-'�tr7S)�O%V@i��,�3a�;�ĺ�S�����rCRGa�klW���$�5~|wY��o���}}��y8wI���P��e���;��o�,�7K�Z:n��D�UZ�Q�ܾ�|*7��1k ���@z�6 �'I���a�3��ˁ�p�0���56���|��	�G��f|�Ώ�3�;���s��}1*�sZ�䦘����rJ����F%��960|Ռ!�.��� \J�wv	��Gq�=B��ڕ��$i%+��#�����N�dR$
���JJ$��g]�?z����)o�����u�ou(&�u�����t��^(M�:���gֶ#��
dW��Cǃ�b��z&�������l���&i�����dɎ2��MQ��//XT�p�7�2�Ka�Q��4_���hblPmCCC����9e���t7��G ������A���;OЋW���X#ڎi�ǧ�J,��_?�V�<�D|�'�����v�x������/��� ��9����B�Gd��O�C��^���İÓ�k./��M<�8��w��yPp��`.��A;]�������dnY�fk�Z���-�tŭ�߻zX���j0;5;;�ے���vʺ�^��Zߘ�Y�e��b�b[���6���;�u�j||���3pq2h���<7%�Z,����籝����~��R�p��(txyŔ��C�j$j(����Q�t���Na�?�|NM���5_��U*:X��@�c�#7����{	�H5��T��������:i�M�����%{<ʒ\RU�a{�0jj)�,�*�^`�^�b�S�	������W�>�P������n���o�?�;5����G��l_�m�[���2��iii9Jf��])�ÈH{�S|ŵL"^�vtKZ����ﾱ�,?z#��揞�V xŗT�Sm1��r�+E���B��I�E�/�[�����.%���QLw����V��g�{�-�>�k ����=���;��^�cit3Ӽv=:j7�[���q��MVK��Q�I����*ݶU�w ��H�G��4�^K�Y �0�]��8J�z�kɪ)��6j�N�Rl�6�5��y曫Uf׿v�L���x6:4��Q��~������P}����Co��<�6~Jg���ĒF���/�?v����|U(K�����2"bʑ׻���cJ<�0!���fl|�+�I?��\rc��?*Fb��q�i8�iY:������q4ug��c �ɛ��g��PSQ���ճ�j������.1*.:J3���H��.�����%S�[�O��p��i�f�U���l\�������� ��p/p��6tHי�+��!F��9hu����x@G�T��ళw�5�� P(]��0�����6_x��XʞN�\V�:aX��|il��3�<}�ҨOyO�ak(K�`6:l�GZR�G3��(`���'q~�/ϰ,X�����n��Z�m��-�F�Cf'��i	��Q���g�����Z��PYM:������o�
a!���Xt%Ҍ�Y�R|
� � \�����D�_� �8�j�N��jt�迟M(!��S���cn�x��T��Y�V[3�[bƗ��R���^&~~����.���n�.��&���Y��ZM�e�q[�&gb�p_�z���{:��l�K�I�g�x_K�?w���4CÈ9LW�غx]��B-t��ז4�)��g��  T�II�@1sX�?�To���Կ�2���cOլ��$��U�&��e=v�5�K>;7H���~*�j��p᪴,n�o� ���w}:��YD(����J��Ƌu��l�*=�lښ�1q��&"��@B�͋�J�2{A KC w���U9�,9�X�$�����,���!���Ð�ȵ;�]��`O#�$�	\��oJ�	Uy����N��G��.�f�P6�GFy%4=>��_ez������E�m��K�KV�d�MnV������E���Ӎ��
��3�]w�:�g��d�Fv���7�d�+A��OfC�DD�z����ĸ� �`�xj�B��v�����H �O�BAv�zd1J�[�Ĉ�0�]�l�~���3F�0�H1��Ԯ���W{v��d�T�
�V�$#�M,,��d��(����lwƐ�*���Z#��������y�4�rؗg�ۣ~u:�۳�y�m]��2�`�z_��Ȃ��r�ni�����7J�Z�t���}����q���#~�z�:V�ʦ+�����3����
j@�c�t�r�o߾537��� R��'Q�Q��?��dLT
�opJV)rY��t����=�K�;ep4_¢C	rz�\���}e����1=u����V�����x͍�<�0j�:HH�D^�BaHj*�����A�r���7:���߶�$7�g��������=�=Ze�:Sy�j���h�s�(9hΣL�gJ��ͣ�K@��K�i���+���IBUm-0� I�<�Uʟ/�~Y�f���c0+�m}�ݵ��h���r��� �bQ���P�`h����&�72�_�6V�~��J�Z.#L������b!	Ck��?��7���T�Cub��ag���<>����Β�_�ڋ�|j;Q%��Q��lN/q��4S�^��������^ ���Z�^�|�H���䐇����	��@���8�����O�@��\1��_�֏7�q�p{�PH7�'����͍�Y�n�l��LF�����+���3�G6���c���#/�(0[���t���nZՊ.�՞@�Ej�Ɔ9	�5=@� p][+[cY>��B3�]����$!Ќ�h10m�1�T�c�OY�@A}�-1������^{+���|�j	���N��w����Qm��{�M��<��c�w�G�����������yCG��J+1%Xv�L�N�6p�����H�����>j��l��I�2P�_l!�G�zz�9u\��������)�r��`K@֪�+T_�$������#H=H��%C666�����*�ХeP�D	�xW��V�f��� }���ng�Y�Dic�8����� $M�x� ������ɂ�{�?�{�M����t�&'U�c:����JS�q�^�O�,x�#��
���h�������C���%�WX�6���{���s�Y�Θ쌊��:i.�ä������NJ$�HtX����q�*��>�NI�����6VH&1d���PRr�CrT�&��U�?5e��D�~#�|lm_�i݊�Z��x�A4�RU6�L��PLe�=M2Е�6]߀:W%e_5���ȼH�L����V�`+�:h�@�ϙ�vZ8�kk�Gal#��D�������.�?�?���� ��gӟ�����
�t�9��_�%1������9kʐ��ߞ��Bm��B����0P@H2�|�,��i��[�?o/�H���P����:��Th_�E*��H��:Gw��������l�
�fl/�c�����W>��~]�v�ӳ��>ߌ�
{���[q�~l�I�՛p�Շ�k�Bov�JP���4� Bh�;MO����������c�($����{D��������oo>���:�����#�1a��r�����M��G���8��`΁�U~|́�lp��)�q?C�cbf�jm-�r�IR5�����u�ad�1%xU���;���>< ���װ�)x�viG�5�P��ȗ��c�S�q����\�t_�_\���9v�9���$��	�7:��?�,�
ݖɍ;��UJF�Nu�](��-��'7{f�ֈ*�uI���yŤ`�c�/]@d�ԭ��[�h(
�ޖ`��`;�Mz�������xL�>z�ߎЭ0Hh>4��~7�qZ
	F������dx����Bm�ea�j��f�#��)�sU�?諔$u�H���py�b��
�ߧ� H���4R�a7�13$�(s���φ<g�;���Ҝi��@��F�·�'G2�K�Ee�aL�Vԫ��q�� 4���e$��ϴz�s?ap��!�&�ρ{�o%*ɗ�ڭ��qli�? 4�}�*�������[#in�9�D��)���n��li�{{0Zځ��s�֋_z��&�	ӟ�Hݲ�*��F��U���0}'�%%W[�y|��gKf�9G�Ht6P��`��{g�z���&75�8�.�H%e5hn�r�f���f�3i(���E�T�BW��#l����?4^�5��l���B��p��n1H<<����p 4���v�"w#0���4�7{>�1{�j���cs'��I�~��*�F�,m�А�Cԙ��u�Xp�C��
���jʓ����T��6xs�X� g�� О�4����X;oP����u~s���`ݲ����^�Y�c��@�y!���GP^�\rXF��B�+C0Ȝ[�)j�|�q/�ە'�%A o���I�g��Y��VU˴�`�%��%.��0ժl2h��P�R����ro�Qo&n�_+�}������U��G~�,����kzv��ȡL�?Ǡ���7�T�v�N�/�����&��j��p�Y�k/�7{�;�R�T�Y�rA��r�pp�Io:Ͼ2:�w���hm���A�BZͻ��a�Y���^_Ћ<-i��]���s{(س`Jn��P�B��~d�[i�Z��P���˞ж���q1���g�c��*gXQ��X�gϤ�2b� ���8�<B^Zp�iQ���4	N�|�5b�2Ijel�W��P҄����3a�hfP�NL�;��{�n"��f�ΤB-PE��V�ދ
��y�X-Y�l���ڎz�]N�7<���v�n�ta�ڃ�5���M+����&\i^,S� ч��`��C�Op����V�b|��7nXuL_���d���;���������_
�}`#������<OH��0�$�u|��$�Ўc��� <`��h��,�is�5��q�#����?��Gm䊊��F���W:Q�^�:[�`B�J�Vw�f�I�ƛJ̋�<W�ͤ�6e�{����{cƸQ��2��|�G��]����h��síp�DsD���ؾ�nw�՞����NZbؖHZ�v�W7&ڙ;wB˴-Tv�8�m�u���-VL&o�g=�":��+Z�
Y��$Q���cF���`=,�$��:_���(;C��%�6Y��B��%-�k�=z�}���~�%̹F�/6� �Z�d�ɬ\��?)O�����A&>u翃�����~D��>��Aƺu~�����ľ�6��e~���v�qJ�r�L�
҂Q؍�G3��`���ц���iK�|K�����w�����_�-��r�v=4��~Ŕg�1C�\j*�|=ެ���~�aB@�q�:�w�!�p��u�����Z1I�0��|q8T*�y!T�>n"��l���Uѷo.�c=F(�s�-�L�[�x����)L5e*��l"A��j���t�QE��ԑ��,�LQ�Ӆ����풆��w�6pn�_���!#"�.y��i�i���Fe/��,L��)�����Zef�a��M��?��$��.�?�p(p8�ej�=�V�t+��+�f�+ �����"�u�`�yM~�/[{��٢�]�^#��6�{�w����c��0JJ	�������qn��.���@}p�L�AV��O�g��4*�Ǿ*�� )9�G[?S���
c��ޯ1�ӨW&{��Z)�D(gH(1r|�(�^�<�����v*��4��j��i�F���\(����t�5��վj���$#�ԋs���@��&��������ٳ$�`N�%�`.Q
�d�VT������/�*�:��-�vۙ��K�f�X�/Gт���d����	 ��glI���uܯ��t���$�����X���r��,����L�4��u3g�kx���Y���57�{%O���@ӵ�W/&�(~���xv{���5<��PH�ۣ���GWA��C�8Ge�k�\C�̂&��v.��L����r�t�*�9<��3T��L��>{)"r	��$((�V9���~�z�P6�|D��菣��/P�12�Hb��T��s;3
�)�Wy]�G*��ٲz�&V��){^��z��g��t��sI��ή��I��V��-29��HN�6Ûq�(,�A���M��)JJր�Z#�H�9ߜ�}�n�IM��y�wc���[���/mWݯ����I����޴���y�vQqN_(i��Z��Y��]�����ۚ�G�D�\f L?Wv&��ɷ!��浉CEƵlW����/��B�:a\��}��D���|S7��0oO�����������B��7���h����V@�xp�;;�Vnۭ3�,--�	�$��:�ٞ�(�ѣ���~q�@�����~��(7�Ǧ?�T��� L�͎%����&;J�F!+�2%��e���LCs��gf�(�a��t�v�^Vgh�����9�MO�:����Pi£��q�m扖�ǳ�ǡ�����S_7�)��l��&r���"z���͆1��de��'5�2������.k�7~�@~7�t����j+5w�x��ߢ��O�lj��!��:eyڧ�7vN&9�ޛ���R����(`q(����D�M��aTk<uT�@�H��U��N�g'[F{@ª.Y���?��QO�Ƭn��gu��3a��r
Ғz�UVB�@��jo�$�l�����#:q,ܡ��+1IM�T��w��sQ�WY�����"䉖��gϤ���ذ�D@q�)�R��)>x�oK��"7$�tR�g㌽�*9�T�̥�����3�����=Ѣ���%K�__J�Go[ۛ���ѻ����N����;濩��sx��U�q�u����o d�d��֦�گ�M�G}eZiBJ�`v�W�*L�|8��\��⨵�������"==]�|���y������"��V�a��_���<��>~{�z%���]�:��%�����}�R�㝂���G�5�������U˴�v��>}J��s~��q����*����[N8����������G������5�ט�����*��š�����_E6��*S֝��8u~�G���#�3�P�y��p5��Ap�8��?Y���
��������z~�2#�"yE�{S}��2�{K�ǲ�������>U�����C�t�D����-a����Ɍ�-�/_>�=L��X-#�ksg���|T�k;L#�ʶ��`����E+2��tt�DO�����(�o
��a}_~�[M�	]��a~" #(��9�s!lޓN��ܝȲ%η-��a撓g2�@���{A4	JP0��r�d�YTՍ�/�����Wd,�o�v��Vzmc#�
�|�츛]П��:����WÏq�7UTx�K�S��?����S��$�I
��@A��h �\Π�!�����?���t�!�A70j���a�w�� ���=�<5�=ts�%Z�ps�wy����F���Z�N�
�^=?�Ӟ��y��m�����Q�iHA�r�<o�q,���7KsZ7&D`5�#]0չ��X;�_X��>��!�TzЋO#O{���d�{�C<w7�1�{*aK;����
�V2p-GY�s~ε��|�f�5Ϙe���=~���&P�ǜ�?�We6�!,W?/C�T�b]�C�h�%*B����-�O}7(#N�i�։�;=�R�ť��hAƀ�J�8����)���4�J�e;�R>�q��?6��)���ӥU0?���,%���O�e)C�.�fE� 4AD���5%�`0�`�=H��P�4F�jҏW���#<??�g��k��1���n"@3O�\3���TPv�hh�7G�2�.��Y�E�`"W�Ö#�'�װ�I�<� ���#?L��5Y�?r��T���u�җ{{�FPi0O�C4fD���ׯ�֟���2/pE�Zu�	-*'��?�
2�VJ߶3��WDA0�U�K5:����c��\���/>��=�a���P�p�)�o?��Xr8>���"Ab��ƾ�_��k��KɃ����N}��o�lm�o=s�`�,���-����L�Z�`��_���Iy��^z÷|9=f9}���8ս�!���a�Z�E&o�7��T�d�W����I������!+8���u
2��?����< VW�g�)��T	��v�פzm��!@U����o��-/@�+��4by��?%<����r��,��N4��jn������P�����~�oi��OA��{����k�k���g$�6�ms���R�#-�I�UZ��۞��=�Lh�B���m��yO=--�3�9�ޡ�Z�c��v��F�=�Y����K	����KBT�y�Ĭi.	D���0ϖqAǭ�g�2~':R�?���T7-�I��D�g	�	�~����m+�W�"�mmvgA���q�6$�Dr��ZA�lj?fE�<�_.	^���u<������
����z�e�Z@�+�mD��#��!u4��`�⒄L��뷁7���7<�,V&����쾇�[N>����l�~�+�urt���U�{�$t��:�ʒ�%�����ր����Jn��`ϰ�e6��w�~�.��pcm�a(���&�t^�_X�0Q��J2�R,f���+M��a��<b0��6wnp�z!ꈣ$#8�]�S��"���8��R���V��!�\�e;??jѻ㡷��=B��I��g�)L�����lYu�ė�Q����C�/!��ȡ��UHŒ�S�WJe�,����:2|Y�-, ����`����^��̞���c<
,�?
�D���g�^�^���w>��T��Oq�9�A���GK&5�i1����-�)��1���� ?w��� ��O�Yjh�0��#Tbej'�ݡ�'��;�|}�uR�l0����dxӵv,Xeraa9��L_�-V�;��m���jIɛ&w;D�/|��q�0�}����P ���[	�7�"W�F�k�-�7�FyW�ΎA.�Bl��ޚ-9P>����H(<�&spӵ��'�bϖ8s���#O�Ќ��Nq�[��O�hW�V"��]�p�p��N:NBd�5�e8���\t���gS�;ю�i�������Be�\��^����=�
�F?�!�9�ۦ�IھO��x!=����d�����M���k.���/q(l(u�hɊ��:'#a��㫎IOt�M��^|lllX��Y�5����Q:x�I?7�d�&����x�/���ux��U��u���\��҇#���qq8�Ӗ��e���G�k��˥��8'*zR�뇒c��}�/��y{��������&Ϲ;�
��y��.�\"�E��7��Kf�й4����2&+0C/�2~���єPB �H�H3����(g��U�![�c�[��M�d��(Zn��s�®�`��q�.�z�N"��&�v��/#
t�rU+�^K]F�o@b���M$���	Y㬀q�\^�N+���\��S+��_7l��`wWg�)�9�+�\f�I?͢�G�=�t�v�dB$���������\777�6s��>-
" �T�5r��}��m���U�������_O�w�5j�英��*�{��i�q�#t��F����8����Mb�I�Yȧz}��K��ѸNO�@-���j�̓M{+z�҅y�a%��Rd�ɤS"O5��t0Q{>(�d?wy����V�Mi��2�C�Ɋ�������v<��J�w�5,E������`��Sw�IF8<�z����`�(0͇}Χ�sf�ϝ�5V��"F��e���F���J�Σ�UJ�@�� �'�$,���[�����Vx��w�=�9	�[�c���CT~/ũ�1���5�3�0%�P���:J(�w{��&j�"��v�����#�L$0R���u���Ojld.��^�Ε���O��&��TU��z�����'�:ϝ����d�o�|�G%��D bV��*������1SOϴ~N��n�p�������-�,[�Jw�6���a��?֯�ă���ɠHp���+2S�XV<$y������FRD���	s��!�HS�"����Ic��<[��ju_Ҽ�b,�m��l��$�W�gk-��S����p����VT�΅ﳧ��ۣM͓��	׫��<I~�Ӎ�z�������Ht��4;7�Tx�S�Œ��3@��.��i����@a``��������-"Ǐ��$�	XS��S�B�߿,֙�TD����,�xTTT���,߳?���������'@ŧ�|�
g�)ڊ"fn�e>�+U�@����Zt���i�	���
��2�>�Z��,�[c5��~����(/����[�6�kƑ�(��2 �����P�5�{���4�����.�XZp��$�Bb!��&E��y��A�1ɗ����1�s>���y+r=�M����O�c�(�F\�P����5vi)���?W���]:5#�_�������d{��@q�#y��J�N��gg��g�EN[l:M�MF�l��ޠ���g/�l���=3gyJ�П2M��`����1X3��6���d�g~�'�,Z��`D"�O��-��J
�5�3�O-�Y�!~�0%��S*�[��o9��O�9��Z����#OO<u|�S�ɨ^L���P���	d��e��Y'1��������XV���IC�m�\�m$�O���SK�!���=!h����i��;'Ȭ��,�=���A` ]����ܡ�s�+d/fޟ�V8��3T��(Z#A��F2ɕ�}��LP��)���jϾ3y��EA4�ÿ!�I|~��}�rX��V4�=��=1Z�>خ�?|��f�f�.��m������Ӏ@�N�.�M7��xAZH56qJ�e��a��MNid�lw~	u�����`�����T5���л��k�И�������_�6< ��p�)�����N{?\o�p�C����� (�o�ě�)I���Qr?V��d1�)kO�qC�>D򥢽]�:`�^�*Xt\'7�2{4r{I�����_[÷�o�#)�#�Rc��!��sl]�Ti�1��_�҄���P�����)����n�sc�|SU����������ܗ�4�	�t�=��"1���m��)�	���l��Q���F?��Fkw���O��O.��pqN�G[O�gm͔���KҪ���Hvσ����Z�Oϩͧ�p~U��_���{��J�Jq2d��~�6��p��@�*���F7�iQ�`ۭA��8[�� r�#Mg4H��@��XѶ>&��>��(�S�ߣ�!(�ku!|��.��k���?�jQ�(�sE��\�]�ׁH��������c("Z���G�G�:q����C��v�����0'p�3kR�LmQy)�u�&}RU�h��)��;X��;2��� �SQa�p�I��l��x���Ã��k��QMM��k�_嶭���r�J>9@�bs�#����n�8��3�xZ���_�>=�����C��Y@���o�\�Ve�X���w65E���}�g@��� K���^�r�\�ZJC~z�O�� -DϞ5@H��K��D�l��\�zX1���&��CG����ƠT��y�޽����{�{���˘������''���>��f������jW�^E�^��˨V�q���,�l�ZM�y��XZZ���
*�
j���c���ݣ(�ds�ztt4�����7��f7X�B�=��h��]k�eo�M��,K��Ǐ���L�|]��0133�ջZ��̙3سgfff��".��ٳ�/i�F%ۇ9SƵk�2���O��(�3g�qN�N�s�ضoߎ��%,,,�ҥK�w�����T*���֭[�s�N�B�lf����)h�q���4C���ܹ�z��z����E\�x̌������:-�8���(�Y}�"�=�!2ײt���2�og(�� ���Y?~�����_<|��J}��F�W�+�2����f�����>f���oI��i!��9�{���"�ipY���������	���s�d��!8���&�A�)~�3/��h��-�f�N,�P�a^3�܀��̏�N]���o�4�}.K�Y�׳��Տ�U��\��n�u>͠2��777�����>������ݻ�W�7C%$I�Y���H!��I��_��������D�·�p}��#_k�~}&��F^����}������m�=�&02�M/x�e��~ԹW���g~�}�/���o��C��D����+��P*M���{��O���i��1��Z�}���ر����������7�[�g�f�9��zx����^�7�ٸ�|w-�� v�����a����Z�M� 6���޿�9ڊ���1���7l��봙~l��4y_�A��ߑ$�����v��ѭr���)���
?��t���?��?�g�<p������o����A��`@�����GSSS۝��)��3�^��0��g�~1�X,n�i}��$x���c�Q������ǯ������2�ES�ibb��U9�@�ݻ�������(S�����Mp�����H�ػD� &"-"Ph�) �Ҹ J�G2�̬ P��-DQ��0H.����:"��RA=�S։�	@���,B*�[f ���v8�Ի��>�vu�F��o���G��ז1�ވ=  |��NXk�*��
�P�I�:�����6#	H� l"�Oi#%Z燄J 3�Ŧ�[!!2V�b�P��Dƈ� B��rf�B�H$![�u��"Rld)�I����zL*�xJ��k���� ���$Pd{�'�Y$��rb��Ɛ1�����K��r�M��dD�0��T��0�a���lL1SpZ/"!bÜ:�ot:SF�<3�|~�K2ݸ[&+6̅_�7:_��^@m")��(�b���2q��`��Doa@K7�d�D4��N&(0C��@��C)��� h�:M�� TJYf�"�Ř6�z$��Dj���B)Cƒe"%�F: e���5�%	��DZ�\E=P�̖�%
z�w�Ek��~�7zI��0zcPD��zgV�:��ט���F�D�fٲm��S[}|���A׉�E��-=���D��d`ź<�@�!�Y1�LzM�"C"J������Y+L$���T�e�$}�D �DqZj#
 �E� J"���A
�b�2E�$ʊ�$�6&k��E�Jk#�Z�Z��*�tq��Y�~E�;���- DQ�,IL�Y$
�c-u���֚����2i����DDʥ�}"
ED($bf H�a��	��Jqgnn��(������9kmh�i��(��ur B�#;:��8���~%t���8ON�(ȋ�    IEND�B`�PK   �R�T��4�� ̻ /   images/7a4be1c8-201b-41f2-b584-263fc50cb409.png 5@ʿ�PNG

   IHDR   �  �   �6.u    IDATxԽ	��Yu�yߚ�r�}����EBb��@		a-�ݞp8��ɡ����glI���'&R��l-F��Q�#�-4��@�M�U�յt-�������~羛�*��7�{��������{��U���}�{_�ԩ����l���4��T=�z�z�V6�fsPI픪�ڨ[�������aj8��<�%C�WYH3��L�9SMG�Ri���f�ުժ3�zs��g+��\�R��&T��ڨҪ���L�Q��Ҩ1���a�T*�7G�Q��^�Z���n%U:ص+5��Qg0u+�v��ەJ�=�>Vz�٫T��`���y&�Ľ?$�Rܫ��`��m�'��*�ʨګ�NoП��*un�~��6�Z���I����Q���0<��})�>}Gejj�z�ʕ��kk�pd�[��[��"��ߵi��Zo�H���N��hX�u��hTvW��.*k��h4����a�oڍ���^T���zke0Z�k�cm���T�w�	t7R�V�T봎z�Z�J���H\���{j �:	ԁE�{��F�{��FN^�Zu�- Vp�Tj5~�|���i��e%p��>>T� �c@�C�*�A�WG�����bP���j�_��{iX�`���~j����x��F��VG�iuu��߹\o�n7���Lw�Ύ��̵F��Ơ=Gc�i�����Jsz�`�U����������Dk�����&g�;v�15�ЀKכ�j���T�����!\[3��i¦������;���t��5V�&��B�2=��15�NM���O�����Tu�h�R�sWj��s�zcNn^�sÁ��)8��mro�a�Z�Vk�Üis�e2�'A@7������N�3��6 �z��[�s����V�z���\�]�f��>~�� s�w�)���uoЫ�S�s2�Z���_c��;����*�Fs؀C4F�zc�6��k4�!�i8Z�v��n�Ќ6���:�X;;Zi_|��}�����/��������XJ�45��ިV���6�٬�F�S�6��f���J�V�;J�]0��h��''����si�֬��>M��Z 3��p��� 5"H��J��̠ޘ�WG3��`��]��<U�զ)�F�:l�氚�Z�GM��`��f��U�pjĔQ{�@=ti�~��&U���`ځ+p�8�
��az͙FO�4K�WKM䓪eҲaeU >I�`�4��z�FY������3�Ju�?\�W{��G��M�f��X{��\��{��'kS��a3��ҠI�6���u�oZ|e���C�����-X�l/[�/Oķ��]S������
�.%ޛ{��Φ�\eX�g#6�A�ҨUa��ҥ�+ w������B�A}Dk�fm4���0�y�c�E�* u�l�0�Z���@�� RL�)��-��n]k�괓J�E�W��C*��_�$�V�V�aT�����h!�9�$�6�j��v��?��� w���?E���fZ�p-�!{y�p��L<��1lT���R��9����r�M�
ʫ�`�HC4�Z����v�ta����w�oH���kmG�ѩv���Yo�#�]IW6��a����� ���F��N6��c��7���ԧfG�ֹ���9+)�흭�;k��;����1�r�G0!8%�Ym4�*���pVEXE �OQ�C���R�	����+��lTk��<��p�f��:,X+��&�n��"������4�w��ۂ`�$�x�^��ʆ�+u80����hyv�mD��0����E�H��/#x�� ;�7��K`�J��^!���br�0��Z�F2�]��z�D�a���0�&[�j����Y$}�[g�MB�K��A/���ty����W�6��W*��0:�����t���:HD34�3���>��O=�p�Ȯ�S�.Y�/��o�#oj�Sn���ߓ�t��P�5��O��޵�C�����J�Ԫ�Ȁ�^���ht��F6�:��4C��e�V��kC�^���:��5��� v������C�3Ih&�;̵�-�A����3Pl	�dɽ�l��M�#�qv7���,��[p��F���r��M��i9�v�E�66�m�#��6Z[[c�Є[2r�;v��]$�t8x�	��
��{�n��h<0^x>͂��0��0�?�Dk���]���Ӡ�{���)�huuuH�Ku�4��~���_�W����'N�Ξ9��c��d��h���2X�IYIk��N�CSb��t����T�I/q�#z��Cw��������_��h��[����la_��;�w�{ߑ�f�A��H���F���:���BlTj �-D�d����RZԨ�F��Ezպ�u�0?P
���f�������.�F��0?j9�J����O�q��Y_�N����ⱚ�:[�;x`v�_�V����0a�ܪ�
H���"+�wSkz:-..�;�#=�� �3V�NT��Fء��I�
�l���1ۆ��W���󎷱?z-����\�k&�����M9 �i��4�X�t��yԅ�M'�5-��6A�477�P#%M��fg[�����]�y��{������p�����7�'����y����f^��[�\<�䯮�;��~�k�O�c�*�s�����X�ô���ܫ;�0�:��۽����qe���X߻w����u��ý{�,>�ܩ����Sw���tfgg�Tp nzj�t{��
7��y�|V�m��F7R��NK�.�Y*k߾}���<� ,*�
�E�"�2�-��faa!���H�A���#�͇\T?�	��r3�*�,4�4��߈�m����І��v�꣙���ph�(à�h�C���7a�1�MY5��u�2� И�������joТ��p������?���Ni��S��m����4]z�4��/_�۰\�4ݬ��w��;��~�׹��gy�	}�������������g����y2�DI��C(+ree%
.����ݯ���}��}�.��f��l���F+k��s(#F0��z����~��=l�رX������,њ�� Y]^Z��߮=�cCr�$ph���6�/--%�.)��f�޽�g�}�fc9x�`ZƟ�p�����ܹsq|�����ŋ^���#G���gϦ={�G��#�M_@{� ��`�]����?���E�f2�tg����>�9#��"�W��vف�-!@��>����"�!:�4^�9Q!�� `HtY�Akz�7M��puZ��ܵ{7��;}����Ϳ�7G?�����t����.S�Fp9�y���0=������>���?����_Fpg`������O?�K���-�kQ8���۲���;�����kp�����9x��={`���3���,�އ~���t(/�o�!�v
Q�"v�ڕ�}�8�ٝ�h����r����4����4`��.����>Ŕ�v6�1�n�׿>=�����o��?w�y*���g�`�xꩧ��wޖ��Xg �ћnJ�^8i7����G�&���ao��栃�V�p��=�W���m� "~|�{�d񮝽�ϲ 7{�tן�0� �\��]��s���}x�]w���;���ѣG;$Q=q��G}t������8��8�����z�M�"�����{ϮԚk}������G��ۯ{]j�^��t�/#�S���z����>�K�.^��馣�Kt�s��j�B=�ēi߁}�[^�����鏮v��ӳ��gN������ޥK�y�w>��cvu�#�IX��r-�V��-�/�|��b��EZi�� 2[���r�95d�L�Yw9�~��J�cCAU������`�28d�-h�X�i^�
�uX��KD�cںf�e*�����z��nܦU@�[.7j�5���6��6��_���Rb��VQ�[nI;w�L�N���߾���<�dT��T?�هv��Ϭf��ި�"�ow������;����=����w_�=\�e����8����깳ggn>zs�Knm%�$h� ·��=��p������1MG�j/_�����n��w r��4	f�&��Hʝ�V���݊ ��qX1���8���V��Vhe�^��[��_��&�h��n(�#���� �n���̣q	�*
���U@l:��4��~,���hܥ���_��w�w�툳 �{y.`6-�ҿv��(6#?>��2/���������7�����������y��O|p�"�yl���B�sp��'Ϟ��sϜ�@$x�?/��{�{~�g���O������瞋nފ��������������nk���c��_������ߊl��y��(�Ĳ�#єQm�)Ǫ&���-�ӿ����b|֘�@ׯ��X!V��a#�b��%����q�Ƹ��Tc:����l@��0W�q�N�\��დ���|�|�y������2L���ް�_c^L˸
Xԇ��(&�7�X��U��1�n���GI�<�.�����;��������MGoZZ\����|������;���LM�^����g�=�tgj��~y��?~ꋏ�N���z�*���E����ﺵ�z�O����B�þ�� �2�I��-o~c�5�������^������G�������w=��*Gsp%g�V���YQ>[9�ґ9u/``um��0[cX+ɊП�N�[�Ƨ�>s��9M�nV;�^@\*���?5�9�y�bi��׼��%�l��ccN�9���ӫ䭼�?Ǒ�e(�3fp�p�����w�$`�����(so7�-Ƽxƻ�g�q@k٨��~��tӠ ��n�ߌ �K��K_:zӡ��˗�����k���	��M�O�����ӎ�����G��󒧯�Uү%�K����;>��_��=���5?7;���G?�?�rכ���W:��M;w.<���C����� �D�$��%�
 $���z(\�
�Yc%Hl�c�������5�m<��e89� 7��U��)r�፿?�m��<����<x�������U^�b|�1�Gc��5u�ž�u7��ny��Ԇ�)�Uw�1�����g���x�
x�*�x7�H+i�/��}~�������2��t�w�qە�;���_�B4`�c�~�4?3��U0'�.V>��z�f��Wi�a�޿���������O��ϷZ�dVpQ��,`�B��H���������������������'��1�{��A[fg�g"�Y��B}bრ�����ejx����������4Rqأ�Bԁ��l��)@�Ӛ&�G蜩�aW�}�j/��a(J 0b���~�j�:[R��<��`��/s�?&��++�V��#��X��/�*%��HK�xU]G��vbJ�Yr�_��~I�r�O&�`0���^�
X��,}�6���dI��(t⦇{$jY�P�u��������0ݬ#�n��}�ˏU>����I~���5�=�w�����~�S��,.�D<�2� #Y����Uf�����[<���kR��o�y_��5����?����(Rn�r@'D����_��Ks�|��;j�c�����7�8�,uX	��% ��X)@�+���\yY�&C�K�Wg���CN�����Q��y�n��a�2��N4O.��l2�
@а�g�cI7�<�7w��	�MIO�(�ʥ��;ؔ�IBoq�9ά,q�D���C�L�8K��w����4������7;m>i��Þ���}�L�g�o����0����'�no����='�y��Lw>����.��_{��������g�x�׈&s����?� p?����++��w�������'�����y�Ϳ�ꠍ��_����ן>}��N���X�`��@�E�簞y�=j<�#����Xw���\}Ϡ7�Z����O�{ En�'�{���`���lq.����'ee�a�'�2>z�e�ў���vYB=��3��%�|�`h@ή���IK&P�wpB1&�L�E.�q1���0�d��g��W�/q|�=�q�:�YTV�ɞX;ELEAU�6p�D���]Y�����S����<����Q�2�W�c5��ݲk��?�t����ľ��o����w���'��?�!&2��(���w}W���~`��٨l�}Ӈ��}�)�i3���2�fP�d������.mԖB�_86�G�XN���/;���P�A���I�ͺ��B"��Ńn���%�|�4�������O�K6��Hs|�'@56 �~Ez����t�LZ@�=��n�_y/�"jDb��-��%������r�x��U�7�ǶE�.��ږ��
�29J����n���t�������߶�4�n�	6�c�(�م{�6p�ʕ<pח����}�o���~�\^^Zt)�\/b�^�-ߜ���w��Fgu�������_��ĉ�Qߔ+s�����11�`ʰ���O��$0� ���GN' �2��
+Ŕ����U�ygu���A�+�4�!E�٘��`�|�?b�*k�
�W���d�1y��q�x��J�Y�J������8X�����U�s�tuf�ysU�����w���iM��l^��0���6��w{��T!�Ὂџ������(��͙Ji-7������|��e���Ѵ!��K˨�w�޷�o���+��4�w�����С���ǿ��}(���]�>�D����8ל�;1�X?����/���3�Tv�H�n)ڕf}Z�GFEۅ-,̏�.���b�5�Ӡ����.J��ݻ\_�ɻ"��H���ߊr�������&k6�Xz�ہ^,��Y7A�����+�Ҏ���ɘu��t���� �"]� ���}.��v�V�˽���b��b�����/å�����"�嵮�&{e񩩼āY��Gx�Ȼ��{.���o;y��#��Ǫ;�8���Ղ�-_<�w���kZ}]�޿��ٛ����g�y���wJ��Ξ;����w������w��?��oy��O5����d�R� KL��<���h��I|�R3��$Ga��G�E���s��n
�r%d`h�J�M�E�֗�5�|en9���qF�!���6�h\d2dp"@� {^��bS7�'�#�JT�{�I"���1�`����C\���O�1���s�{���|�� ���/�mҮ�+~7A�q�W�"��|��޽"<ޭO�C�}|V�)�ehEty���w�yw����ؘ�����g^���zh^�"��lk��YY�y�7_�׾���������F�y�OY�������Cϝ~�飿��qЁ�3R��<�����Rg=D��st��e[����	B%v���<������>�G(�"j����e���d������g7���䃻`�ar#��E~4���@w��2��JQ� d<g0�-�ρ�/��ǱN��8�چln��R���pԜFx��4�^�I��\�&�9�����HW�޻i��՟���=�����{ｕ���ﺀ]����Y�� tn6�'�X\h!|𶩩�S++�U�k�d�k��>-���ɓ3-�E��D�������z��������/}�ᣮah�X���y��Ƅ��
5�ᓐ�� ��V��4VeT1a�G�t;rǜ?���9����@��(���������E�aۭk���b�Կ~l�=��v"g&M8u����4/��bW�ѳ�+�l�ٕ���:rJ��\6�|݆[��tH�+N�����Xp��"���r/f�k����t�_���!(�e/H�ۻ9��eC׉u�]�|W㰔������ df��=����Աc���_S�?u0�8�o>x��W5��D7l���<��{�a�"9�v�J�����0\9��c���W��ڣ���k7�v�.����]2����\h3�ef�AD�W�#L��o��]��sy7�b���m��e�X��\�l3��Ï���h��ޏ�j��6��d͉�[�R�\b��a�n��Xg��Bf2Y3M�`�x�����^N����`Jy�t<G[ۇ�m?湔���Ky6��>dx�    IDAT����O�O�9�g{݋�ڌ×1j���R̱�l��+^�џ�ٟ�\��$�&�1ק����=w���똼��:�����W�ugs�{#�i���TR�Jܷwwj�����4`E��e�Q�VY�In`u0qiy)Ů�̳6�-�6�☉'A� �LC3I��.�6���~��C�IT�n�aC<b����iw�x}~��cr.{1�bm:|���74h<�Įw�ʺ���/������n#f�����8^8.��z�N�Ӣ��nᪧ��t�t+�%��I�W���,�Q�z/����d���nw�L��/]��L�!q�s�������_��_�x��_�rՠ3���?v�-�^�to&��'�����2�|m{�����-Dk�klXJ�����+��8nip�����T� /�AN/Q���bO��s+���*��ƈ�5��P9�w��9̤=��dw�KT/�-�4�	�{����i�VByqe���p�W�yg��W��{Y�Ȋ76$�̬�(*o
Q%��Μ��7�]YM��N�>�����p:��P��v����ŝ�m�̯9t֞V~_�g�,��4�[�b���~��~f�~|.�x��~�]���2:{��`���`��UR�w���f��;�>y�q������c�f��?���7��9��G�E�<7�����'��X�����o��'�!���*k�i �6��c3QM ����	�D��A|OЍ�F�FL��_؃�,=!/�z��	b0�?f���d��U��\N�;���r�V��_H?��ߛ~�'�}oL��c���z���;̬�7�k�c-Hħƀ�=������ ڣ������}��!�O1x2=�!��ɁhЇ2+��eؽ��$�^�[�z�Aclo����x��ڞ����a}��ƫ�gY]Ӯ��/}	���i�'�|<T�kk����;23?�.����<\����]o֏*7�(�����G�{�P�͝;{nJ���-��#[��V�пkC�ɀ�Z�����G� ��8஀1TS������?�j"B�����B�i)\<89y��D�=s�R�;?�w�;�y���׼P#J�Y�ȅĤ{lx޽�^0s�e�+�9�!�� ����g��w����w��~��>Ė�+�j6����l��W��(�n�4/��!�F�I��<��:�=���%�k�Z��-'Wl{�G�?���c?�c��[oM��ǂ���vгէ�կf���3�v^Y]�ET����l����uZ��ڕ��Ȓ"c��F�u��r@��a(Q�~՝�0�;�t�W�� 0:jE���c<2���8gH#��Dp�<K���A8�$�O����Jٻkw�����t{#�G~$���X^�H+4R1M�⍃C�:K	f)o�%Ͻ�3"�u��"����^��q���tӾ�閃G�/$;�u�?'��^B�xH(�$G�Ř�k�'���k�y1�M�1��{2~�帓F;/M���cq/~��]	�B`��Jw��#I���ߟ~�~ ����+1�T{��T����g������6�iHC��NW�?ɔg3r<Qj��խ��͹ʩv?�yӖ��% h�W#s�1]"��ݳ����,U��W�^���{L�D0DD�=B7q}6G�ʂ{�?�?�~��~*zOv�ݧ�v +�LM�R��@����Js	��"�2�6lv�Μ���"+�s�3gӷ����w���c���
�|N�=݆��5.e�T���z��I0Y�k�O{��)�-���Hw2|<�G�>���/�|�L��Qc&�����Z�݀����/~1@���iP�_`�Zm���5��=!ou&� �W�;v�sG����÷m�3���򣜫�&EZlp��^F+�xg3� ���\B����! �HA��n��wWgi���Nd�96�J%�F,s%=t�6��\�cu"�I?��ޟ~��ޛ��?�����/_f��q�+�zZ\��a���B�O�G�xfc3皱�� 8�"��9!:��Q�NU@�8~2���#���ߖV�	.^^IQ�'ϞN�◝bI�;z�Ln��c�y/d<���=�ԡ�6(��*NbB�����qz"bO�����u`Ᾱ���tB\���w"cP�d��;�U�+��w>Bw�"ꓞ�Cb6����=�G�%�%r�jS��^P|� u���<�ݿ'�20�ڷ� ���$�z���` ��\S���[V���o�;j����ڿH���:�I�R�ܙ]��}+�פ���yw��Jq$.�U;�ڈ
;w��xn֚�s�A�_~�{g��U�6�)I�R�ڳsGZ�t�6��e�2���X��(��UQ������:*�U� �� ��,�an�R�f{˂�m�4���������|:�z�5&�R����r[Ȣrw��L�������	Ĵ%Mt���k�->mi5IG���V�H�Bs�͠��`�r��d\���	46ƥ1L�d4e�=�=��=�Ju�s��&���m�~���PGG���y�Ec��f�v�S
�I 춞3���eoȫM�G�$V�&��zZW��9U�l'�G��V��8 �ҕ����X����t�]w�!.'\z���1���HZ,ɽ�]��}�|ZcAm�6;]��dznW�8B}�͙M1E��M
�9T;fgL���F+����3�G�T������ԌϞ9�����Jg�.�U�p��.���E��Z��^��T��aB=WU҈H6���Y�A�U����M�n�=ד�'S(�W0@j�$�����'�o���GJ�(Ø�n�5|��a}�4iykLt��aG���I�Q�jm�ڵn�y���w��<qb�I�>0�=��9s�|�BX�R��,h,dl�3���E��eL��;�
�L����g�� -&�bU'�._:����7�����I���� �9��tGD�H���u���@�����_XS/�����`F$k�����W�퍛I��`�TnL�s�q�Ip�*�g��K�2х�2��uy��w��">�ܩ�O2=�����w�5�K��w�#��W8����$"4�<�cj!��wa�a��H�B��,�|�n��:-�wK_��R�M����\��/�3�-v�UZ�=D4p�h�Vf.���Vޑ����y���>��K�R~������!���tkz�aW��Pg����=��gb���(�<o~b0�����j�R�%�<��X���D*B���kz�h���5�񹲲�J����p�}1Y�L��ƨ�Ђ �yuWN�J��Ҁ��2;��h:jk�����BL�BC�1�x=��"��R�yP�i�Gn�����?�D:�[ED��Ag���e1�-1�D$ٍ۱W�*��N�G���O=\���Sy�M�u�政PQJ�lț��!�Rli�I �n�+\�pk���1Lwm=:�)��T� ;��~�?��������Z�-�:�;��z�'�2C�G�՞��*`ɉ^����MfGjC���AFs3��啥E�I�:��p�(�8�n��c��[�i1�.s��	���Y�m���]{�&�𨁟�'�8�y���3'�4@�Xe��3�	Q{p�S� ���p���rڀc;Pu�X���Ȼ튬��iT�jGPq�/�_�#}B���A��H��M��80���{<A�u ,�bn@���6��t+{뷥{�}]�(�?{�f7���W�*���X׫�0��b�i|[�վ�Rҭ�W�:��\W����D�J�"�M������K��p�˭����^6��uc����/|�~���[���Y{��z�F7?����}3d�A
Q��N��~&���	Q�0�K\>oAo\�lY���� ���� p���q;vK����u>~6��}�8_h�S�{��kp͓�}9�/�O�����Ѭ4��S,5��0�߿l����"�Q��C�'r���54B�;������!_ I����J#08�>��	����[̊�h;쭧=��|���6�z�p�̗K�?��\&����'�oV֖kKK7c��xs&cis�r��������f��>�V��h�]x��lH9��0d4�g������jL1R�J.$sבu��n���+`s��a�x��~��ʕ��F|pe����& �#�k��HX�( Vރh�W��W�L�+��ь镟����M˖�@<+����-oyK�G?���Y��h0BW>�\�s/q~�n&d�?�h���Ӊ�T'�,��ڼ�m�В�9�ީq�lҩ���
RW�y<G��$.E�S��&NդV��ĭ1S�R����O�?�h|���f9.Ã��hI8c�m�i7~j����sHP4I�u40�� �T��Jm�"����(�zy7/ l�.�:�9�W4�q�e+�\���S��ǖ�]{����)y�.>���������ǉ�����upnN���8g���ݜ�\�6��w٧�n�L[����֮�*;�LI{Av�w"�,��rU��6n������/��ϥ{�]/,q$�M)k<��G�F����s���=��� j����i��5w9��	`��\UY�� 22 gZ+��(|X&]D>_ر��E�@�Z�/rT������6��a�3����~�i�H�k⦶D �)�f}*��*��`2�f6�~������v� �RS�C�y�x�\C�vG#}��u��*���>y�Y���2)�j|πͽ�n��g�Xb❚��d!DF���j���l���zm��޽/����p89����B4S��� �%[���}�p�K*-��׮�+�˰7/�{m7�I�����ݖ��?��t�+_��,���C$oʦ;��,8O<�x:�g��9 �gQ���"(׈���@jED��8���LZ�f)�x�7'��a�e_h@�sH�N���K����N���,	�R>������"+�X�AW^������&J����Pi��/|�ߗd"��R��_��y�nU�t� o�{a�����T"_姸��r��^6�F�g��Y�g����n�\e��:S���1���Tk��Ũ�77̹I4F>N�68T�c����f�hip�b��d��f�6	q�FX���X�r	�sӄ�$����3Ǖ��>7�/?��;����'�����4`���g>��t��ϥ#�ȧ \zp� �8]8��r�=��gʕ��I''@�4S�3i�!�Ѐ�j3<yG�H���x�w��~=f�؁���j��`�\@eAN���~6q-M�M��V���6�r���}u,�������S'��+i`K�]���+!��%<����h�lD�VSh�s�؇�Q,�N�r{����f���
'��	����c6s�����ZҎ7A�r�oݪ��O��i�I��������	�L�=E�F͹p���%�����N`1&�x/�;
[(6�/a����7���W[;���E���ۿN����L�?���S��B.?��G����t�-��>��5��2��2mL% ��Tī�Ь�����9����W���'Ʋv��!��@`��9dcW����s|�δ�N#
]^B� �X�iL��-∹�>@����w���ѵ/�:s�1��-]F��F�~�s�Y/=|�Lڳ{1-!�HJ���1����y��VM�4�7	�C�E�V$�ա��2�<gcrح:,75'��lk�,�|�Dw��k���-Y���͎z����ʿ���d�hV���lo���+�-�o�/��F�c. �Lɸ">?V��3C�iL�#�m@?��M?�C�M�;L��Չ����i�w�s�O����i��*�r����. c�%��D�wbG�yԡ�"�X.��+1o ��/���j���������i���YH�j4�MT���Sس��R�B1��Qp�<1p��Qıspp�z	�3�����T��5*D,�^f�ٻ��c�_����Ef3�\[?g�P�c�1�1C�\��ľ��۲��M�1L~.�.I4�N��l��ڵ1E<5�ůq��G����{`�C؞�tN+���$εK1��K� ��(���k��ߟE\q��#�b6[,��b_�`���Z��7i��~�p�U\z�ь���Mm�N�;HSgܡ�����N����ʙ3�>=Bg�d̀uʳ�q�i	hMɓ���zS�U�,����q�v��k��^͛�tz����QE>�.�.l��ľ�H3`Q�"��*.�Jaa�M��ʙ�
Ո��t�|�5�m��ťt������ߙ�Yܛ�<r�5�q/4Y�I�����?�5��+3�l������L��Y23a�~\�>��\dKT�M#���ڨ����67Ĺ�҉v8� �����n���Y->��(��>s��-Ԥ)n4>�4�� ����0�%���~>�t�p���^���Tn����G�U{?Y���-��3[F��"('W�l?��ט�9���rN���s�1p�B�p��` �<i95�;��B�^j�A����q���!�Uq(��^e]>��i��KT��� Xڅ�S�|��o8v';�6��J��%�|��T6�7��,�VM��\�d�����~� >ק���a\�<WX�Ӵħ�/��m���eE�YcsL�5���������?7���m�Enؽ�~5��8�&" ��J��M.�*2lzɅ��AhʩT�7���F�NNeoFăa�f�n�@�'���P�~:��fn{晧ө��J�3s���I��#���Zѥ"��GT�@�2�������L�Ϧ�Y�vd�M
G^qs�߽��*��U�ˈY�d b�3�ӽŠ�M�tÔ8�y�&\U]e���j�(0vP8B���&~^�� ���ͺL���W��N���/=��	��ӈ6�g{/�Z�����b��t/��=ב�����rz�����l�+zD���
Ӳ�S�]���W���b��;�!c�{>�__k�EEO/W�\U\2kf�e>A8V���2��(ﮃƖ��N����*L�G��7����w����ҿ���v��B��b" �Z����@����'���� ��}�tϤ���d��3rx�o�L�z��f߽L�����=%ki�u�s�u������v���3�P��5�c5~�͌'J�@���%�p)�K>�<b���P�9�P��O���#�D,�4n��Aj��F���M�N ;s<�lV�[�I�?��t.�L�-�l��w�˜��ft�0�
=H��g��!����uFP��ɍ���a�Ϟ%4Y�ųV��?��`Q�GYۺ6�b���qbt"�"T(�.̥%���Oͽi	w���`���;���N��i���S�=Ϻ�`,Pf��:O>�>	t߷9��'*����W/z����7|����A'gg�d3L�4���~�QA~�T5��hE�Z�l�K�fĢ����@� NTI�/F\\:#W�n#[��3��ʠ�"{�wltJ���U���Ï�8�3����U�i
=:/َE�tZ�U ����
����N�O���34�@q�=ߔ�L�����ʈ�#l�� {'��C�S��̩��t6O�6��y�V������.PK�J��ٲ˸���|���.N��=}�u�d��"�<C8��Z��&s-��[\Yq�w�x0{�6<�Z�@�]�f�f��]Fk��
��	]�m�]n�z��1�,w������OR9p*����,�b� o0�|���=�;p�.�dЦ!8�)Q��)6 L���C�|>b�h*��;�B7:�1cRn�������\��o�����E>S:m5/gS��
m��(�zQ��I״����u�������\���KM��Px�
ǐ��S�<�q�ƫ���
�����q��C��;��bV���4v{F��R��5X�jg=�+���."����L��r�}�X�\e���n��]cʸK�]$5@��š��jYu7Y���R�R�r/��%�f�m�>�+W ���=�r���MG�
��	4'J�\��~ .@ѿkܨ�    IDAT���i/����f��mqn	SM'0<Mν0�p��#��=ߛ���J���Ui{Ӳ���XcA7�E��Efo3�ƅ�U�+����_ ~�����ao�r~�rN��ڕI�2@��8��q��q]9]YhTl,�o~�I)z�3�E_d���wߓ承Όh����d<�-딾�6���178���D4r�|�-��U���<b	{�5�nK�N��l޽̓v�b����5+��^�ܨX�]-��a�[e�-	�ƭ��~/*���[�R���{)p���_q+���XKN����^�'���o���1��0�OV>��͌��O=�N��ob���$)���h&_������U�jw��n��hɩ����+�Nm@���3�ɘ��)�A��6VH��^f�+õ]�!'W���$�w�1�֘K#���2�&�!wg.�o�3po��Y�z��'�����xi~��4˦��L�_�1`><��^{���矤�6~~�K���.�BN�L˘��xъ�d� �ԅ��f��8���+������ɺ7��.ǖSkWw�;��6���Ԗ��D��~C��ر���#id#�6�9Y{N�'��{K&M�dz �1�^�5ig/My.�aIr��؁\iW�!�����RbwP��S&����g�MSI~�#��QA��=!��q�������m�#P$N�Lm(������Sl�=�� ���Ɣ;u� �ˠ���U��C�W~ﱟ��������ܝ�e�<�P�-]A Y���"��&�ɷP+���;M!&bG���=�qc?P��2a48^x�D�P�o���txa=jG��a�̆�T���sQ��2`�N�q��y���K�}�2��W��O^�_	��������ۚ��wم������8�?�����(�ҋ�=7_f����R��B������l���}�oy�C��v}���l���O���#S.�f�?�m�e���4�� �%����If�����ʼ��Mk~G�^D�/�ٟ��>�.��\�*�ԔAϔj�n�@�*�#E��T�2wpb9�y֓�+8�j�dE�X.�xY�(�BKa�pC���Zk%��(�Lr:ζ�]�p�=;XW���f�:y���M	���8h\j8�7i/�=f�x�fo��8�sWUɻ&��{�����.#�\۸��4�����)�L��h�֎��Zn�!p�l�'S7
�Ի��:�9v��NrҘQ��/�.s�ܽ��hW�OƱ��mGV�'4�wя��w�}�S]�+ru��C=�?��8B͡�jЭ:(� �xT�~��$�3�. ���qR��1f8�!ו��d4ʣlh�T��+L�;Hko��i8#���j��ĲE%�3�̣?�%� �q�+ ��0į�t��v���� O�K\} ����9�P�^��Vqe'�ܱ�{�|��dH˝E�d҃6���U�d}�z�S�c�N�{�a�W]w�uJ\%�r�wq3�Ԟj��y���/�����ùy����t�����z��*�n�*א�Z�Gf�D�ϚRHߣ°�^�����8TMł|
mcz���S�����T
bXy:��3ibՐU��7���չ��9�6N�i�Z���No�����t��'B���n����y�yF�����}w��	�yf��W�bBrC��(�o6\Z�'�hq����co�p��+󦆈(�D6 O��!�=#���{���m>�t�Y��(���i�<�� NZ�,���A�;�O���[��R��;9n��Wȡv�G�bL��u��8}�2{_�TH�D@�t�*��ue�Pyө�h�X����(N�8����yAQ)LT~T[k�*�gk���q2��O���3������[n��@�XR�Î2�X
y�O?�R.@8��E�-��AbG��C���x���)v��%���W�F�md� ���K�|�
p�B8��8�3i�r��q�J�ҋ���#�4��Q����[����Z�ӈ�x����Mhd��?����+���0�<ɦ�U����(�)���:$��ȏ�Q����u�яW�� ���=�O�(G��+J\���ɸ��H�qVj=�zis]�
~��۴V�YJ�ϨߺbH9>���_MJAlW7���3��~�Ζ�&�.ݾǃjv�)`�~�Lz�G�h�w坲���A��KP� we���ݜvt�7����<��vz򋏲����&q�%�6��sPF�!V�8v��3셸���+��	d��gG��R�B�ɻ���+U��
�bo|qR-���v�� ::ɶ� �Nt��=�$���%ݼ�u�g�2~�C�׏��&M	/(5Qd�1mC�~z%���{�k#�VIbh��p��:f+��x��f�Ih�A8�'�9
2x����������)v����ɰ�LBU��_f�ȑ���E'\ �����I�����,ge1]n�*�Q@T �qHe�D�ͺNd��G�Y��H5MsN�i��C���ś��k�J(rDu�+;Fz�l/�&x�[���?�w��4��,4 E����e{�6M���8{�	T�zu�*�m�r�+jq����|������E�j�L"�@�ٴK}�Qy�*�͌l=�>�g����WBL��^Ϯ����r�R�L�,%�W�o܂
}>E^�.7`?���[\!BI�d�B�����ݏv��a���h��]������7��8�	9��+������	&Ťj75%�H���{A�I�@���7Ϡ]`�b�"�hQņ6�M�R�Fg���@�b�������`	-X�["M$8�)�[`Ƞ7�2��F%�n�c�θQ����A"�� �Ac�}��ZCd��|���сY^��!�A�n� ��]7�� ���36Je�h6����z+�.T
wk_��ʢO��('i��1�s(�)>Ðf]�y=s��~�=;��9	1��X�&�٬�<f�
��@)�ϥ �7�cEL\ž�_�o�n�������@A���'O�8-�t��2�3s�>�E�4M]�i���Y���M�z��SMO>�t�Ϟ>�P�f"��RY���x���&rӍro1��\�F'MN;7� ֍�5ʝ��"Ϥ3�ڦ'���lM�ȹ�(u$��l��=��g��L�jLu�'�vլ��x���I�����{ɧ�r?��8���S�;�u2J���<�q]�7��b�t���H�'�+�fƶ�k&	2��]��-�𺖮��4ۤ�=����Τ�#�xq�;֕o��x�=�-�w����dAg��\�[�qڻ_��G�\.�'=���9��p`��,����w��`����+�W�.Wu@�ϨP<x�X�b��B?�!BO�#��QN�J����G?��~MŸE�Cq��&��D�2��L�g.��g�2׭��ix��q��ٸ�Ճy�e�b&ӑQ���ʻ���&o�,��4��-�]�����s�K&<��%�.I���xŋ�����B���|-w��3y�21z�Ç�~���1 ���c��r3Ƶ_8��L�Å��L�Z`X�r)�LS������t��[�Y��i�W��C�"F�(s �J�y0�B�(�؟v��i��'hS�Z�O2������[���mc�!D1�SS|q�w?N�#Q����3��iq	h/M��~J����h���̻v���8�S���W~j�u��y�Q��_�l��K�����{��vB��$K���Ff\BJ��Ѭ�v����K��5o����X�IfA�0��|��f����"m�n�Ҡ��[�J���p�&�$�Y7=��
ʪ��q�XQA�l��G^%)��>�-v쬥�_z(�X��]:��z�xUM�渂4�p!�#�嬔��6Ċ�A�jZ�4Uo�Y�O�sY6�:rw��=hå!����ʹ����@��>c׃��6�lE��{���:*�
c�a�^�	�9D��ǭ��_�Xb��K��]��3��Lk�x��@{JFLs��}��ֱ�ԛϹ�sc-X�R�/�R��N�?�u+N<��g�&r<�vֹ�mϼlK^�����N�WBc�w�62j�hJ�-���\���G~���}ҭ<O��l�eiL��FQ��4kN8/�]��1�c#�1�/?O��t���i��<j\�R�h2�v'+ *�4K�@U�+ؼ������!�G��4J��g�n�z�q��R��U��v�<>?���+V���9�Uęqן4*�+qz/v�^�,�O�'�M>?��G��%.�Q�CQ�Q��/�3�/�z�t�}�;uO9�6�ġ<%�ϓD(�*�(�X���(�fl���e}�\�V�����g%�� ��p6.�C�W���
�\H{�:6���MԂb���v���"�U�g��B
7�3����@�d�GZH !y����R�Є8�2���3%�!�O�9->��`�N��<�Xā��YW����yv�	�0׵�W)W�Ǧ=R�Z�-��{�W�y/n>;�_�.�O���ne$rx&�#/�!=��I#J�fs��4�Z�&:mz�8*p�E=��@�%��^�}�c������]����ɾ��5����D�I, ��#8 T�[��\2�C��U#P �Z�k/ZR40eU��h��2ĄqE(�X���E<%�F_��x�x�L�d�Ы���d�S��]���n�vW�C��(��9zzo��~Eg�����2n����~�5�=�~J~���v֭��g�d�ʵ��Թ�'*m2��g9��lj��Y�s�(5�?���E��yL�YcQS
��@P��F,�o�9��x�	�C9�D`XeȲVqAbL�.�<P���]�'D��j���,� ��͑����R]d
~N�8qt�o�T�m��z�9�oEY���%��(�"å⧔�<���W�6�I��T���\�Phf�qEx~�mO�/h.s	�t�Q�{��'Aܹ��Uc�d��uoyʏƭ[��0���I�4��F����e�kv�<����S�7�ڼRn,C��	�~KW:�S{dC(��t"%�T��&ʜ�qb_�Ѹ�LF�+���h�o� �#2f����rq3���+��	ϓ�RI�ʗn�s;Si�jI���q��(�nu�+��X"1'�c�]��EOd��7��A��`l��Y������]��w��E��2/�[�?y��ڦ�ơ�v��1"�q�tӽ�*<��n"N�1;E-�{�߲K75.�r�jQ?����f6B\RtAl1я�c4a��U)��%���տQV%\�7o�\��f�����c3�R�=3��Ʋ��2fHp���)�'��䙕XfH���R���R
:i��/�p�$������6�-Q)V�1&�D�'��g��j>W��K��	���p\p�yw٨������o�ek�vW�ɉ��+���p�r9�x4K^�Lp+�N��`΍"�&�"�d�uW����ރ��1��z�HO����!��qk�	c�^I�k�盎Jw�~�xL�'�[��l���0�r/>�~��-��>J|宨��l����E�my�#g�q,_B���͡�zy&q.^�Wa���5qN��۵#y2�y(��n�BD�����$����s&^8dhS�Icr_-����0���?z0*P��&�<��6tYk|�����qؕ:�r��KC�S֨�膛���>��<ΨQI�B��ڱ��S��l �4��%F���b�Ʃl,��g��J�n����2ZO���h,�߸������r��.u�����LXIE�F�S�(�n�n���a&�e:y|�{ae��Ϙ����ɸ8�v�<;׵��Fݵ|\���1�v�og�x�-�x�s҄;)�ٳ'�c�� pe��1�Uc��Ӕ�o'�����f� ���`[��J	VTLTkT�r���k˱8^l�{�c\�]N��ӓé9�r�J�AZY��G��e�h��Rc�wcn�*����Ԃ9-t�Ư~z@���v���;�?Շ�P������B�E�z�7�(��vY6��Ǹ��W�uP��H�OmH��6Fp��H����#=�W�����L3�DC�ԏ��|E��3	҉�!��`����ə�তY֠h��ˈL�׆ g�i��ш�ǽ������2"ש_0s��
�\��K�� aͤ�)�;���`���@.v�U����Le�sL���@	剪����̠����$;P�Ո�Y�sx|� ���\�P�� p�X"J�h������i������8g���y��L�7���J�of)0DY�Cɿ�&i1pl K�B�w�!�(�b�8C�i��pDilҧ����|����>f68�\��p�ݒw��c�����9iv��RZa��	m<���G��,�-
P���^;�K1�/X'�v%���Y{3i7N�d\bi��h4�hM���ű��:�x &m��+�p{�neuu%�bJ>����	��Fؖ��Z/��LU?�g�}\�ؗ����m�!�nN�>w߁�|��I
�u��:��YGD`됭R4��д�]���SE��w��;�O�[P�p��nK~��}��1΄N����qܑ��,��	=6b�x��g!���UQ��'	�f̥3��⢖���\���a�aXXa\�H]�A��p^փGħ_�/�(�s�l�L^A���.^����RA;Mq�~�X3!�ذc�!�)X��?�ȱ�<F�+�̤�g���p���V�/�$� K���终%C�s賶#87*�ؕI3 '�[]O������I0�]�+[���C������G�����x���_F"�
� �0c�����G���Blh;��-� qҳ���=�����5�N��'��ES�`ײ�c�{�A^�:=�B|\�5�S�0���p�&��|:\�v!�s�3����)��p6erS�1�H� ġ��nQf�!)�`l��z��(�,�xx|��S�߯/(R�µ�XS6�n!������A����+~J��x,"�'��/��ӂ#���}��K�G}.G�H�գ}87;�)�{ �
rni��`8����%��g�-��z��3L�|���a��sQ�\�xMO�H��̉�-��^����'3���p�9 %7�3�pSzF��4z�~�<�A�nPX9u&��.��l`��j�@ˣx�g��вxn���ß"_�>*�Ԇ��C|�Sк����Qoƣ(1C|��u�)�'����7@������Lm��1��8��J��K�r�i`jn6�O&$Ի�i+�L@�,n�v��i:�& �d�{�cm��x˞����e?9�����g�A�Ϻ�@BQ3 �/������p�h��c�w������")��绗 ���,8�-
o׶�X`�)���Y��׏�������A0h2��!���Y�	��� ۅG~�`�])}�y�*f�#4���8��1d� .#j���\�p� Gu#&8yU#�D�i��DB�H��� �
j9���*���y,��	�d��%�=ӌؑ@��ir��5�=K4�.�q�����c��F�#����{D��+E��ORc����3��o�K}�z`��`�4��LS�h�[��؟��s�My@Qư��g�[i�c��٨���e���$uɚ�{8jJ����%z�Bܒ�R3�cEX +�g)�	'󿆑c�0� sx�k)g�S��$՛o:���
�?�#~����Ө�:��z���tQ��N�ʋ�o�y�ݐ{Q�O%|(��c��` �,�5N�m*�S�~y,����3��Ď�U������~�2��թ}t�Iy�U��#��q�3;�1c��^�g� rA?����� ��0?��'B��':&�G�6kh�t�0��]f���$�H>����q���"�[v���u�U=��&�e����˰d�A;�牯>�2�vݥ%����"��}Sv�t_�OM�%�L���'K�5��w+�L^�X�r��ͻ��n~\���J�RQEbԘ�ڷo_�}���@�.��AX������d��;wO�m��]�\C$�4�s���'RJ�,�*-���=~+�ˏ>��'��)�Ӟ�F�6by	}8eS5����9�(�    IDATw�3=�g��&�Hs���<��_����3ir
GV���7N��UN/ӿ�C��(��ʹK^J����[�_{�7�����n	v
�W�c�m�9�_�hO3�6jN���#2!�q	�`��+b�@.��O"L3o[�B�)���R�Cę������#�.���^@>t�P�g��X���ඞ�z�Uw���>�X���'��/��Q�H�/��a0�"�n�A�z�mX~?�md����yn�K�e�93{����_��:�uv��=�:gyZpw����؞ECq�˜'q�)����g{����ۡ	�Z�GS��:�I:ƹ�p��F'�e���i�o�_|��#t�-NЪRF�J*i�g������J�/�I/��-��ͷ�~,���y0B ��C޶��+�(^Z�>��Y�ʍԼZ��ze���jYT��$��4�����9
O�̈P�s�Y�sC�~��^�P��ٻ�@����Tf!l��R6��@�ZF�P��R��w�h��IS8�r���zF࣏>�n~ű���*i��c-Lϡ��0Ts{w�[o�5�<�t�G�n�A��g��t��G:��G�t�a$�XDðB��k '8��j9 7�7ה�ʳ�=�S���F��i�:�*c�4͢,�Că��Q�Vz�b� �F�=��ic�*^cORz�V=U���t����;�ǂ$ft9��A����Ȅ�~�a�'�H$) �?�j����r��ز͜����Z�-�\��S���������W�rD�K������;W,�hz���+�LX:U�Uo1��P�̖�����{d��ƻ��2�	O7�lt�����Ox����/����BT,q�T��c޹/���4�§�l8���НU�!~bC�+�j��˙U�
��a p��/�l���,W�ָ�+� 	��PM���Xbu��&�'�gt�ɱ�VΖ���xl3����"�q-��	&��l���uΰ{�cS�Q��똿�Ӿ���F~��Qz��7���z�g� [���sg�rZ.e�.�Y���N{	 ��)륷��>s�Ro%�ڗ��]�^�n�z�X��b�b20�ʄ�E�����z�O=�A�!s�9����pfpi�@�Հ�� r�$7R����R
�]�܅�Q��Ʈ��%pa?w�8��[_�^`}����St�뜫� ����S�Z��=��9k������V�!%%�Fqj�-_�����p:}�SL߻@}�]�b��{�Zŝ��nڵ��q�B^']Lp�@�h˕,p�q�N�t�dތ��l �F�jԸ˲��1`<N��Q[.ӀOP�5��(*M�Dx���#�O�n�o�W�iO�U�K}��2h����F&�FFw�C-��u�������;�b���9�u�1`0��L��>�	�(�d�{y��h{hݳ����y~�zS�zU��sW�����HcG5& *��W���b\K$�J4ѨK"*�(��Lڤ����z��_U�y���y���߹߻��۩s��;��>��ϔ6�����d�}
���H���A��>�����X��`�Z���_D�}�fX�dr��#�0���+}���"�2H�hL�K���Y�u,��!F��ƕ����h@�_�}P'���|GrV�K�}/����:c��r�" ?OZ�Y�BP���R����o��%�o>�!���Am�� /}��.�ZX�ݺ;�a��G,����h�*>��(6�+;#/mCf���F�]��9X�!u�0�ԃf�*�W�];@��s8�B�-�����'���L��P<� ��my��`�[�Y���m%U��.�\ i>�я�?�]"��$劣㉇���'��/{�|�?}�����*�ts*u�G��&�,�`25��s�	�GZ^M'Ւ�P/�Yw�<n���*3x�3HK�GX rP��fGل���byy�C�� �>__��`���Y� �#dx�0�ut�����:�A����*Y!�{�=Y�ztB��]�=|�X���B�xɅ/��0ccՃp'K�z����k�{�A���6ôv�i�a�̕Z�T)�Ç���¾(�[^�)����ujXǛ�!
���������~�BwM�n�Z7%/�ҕ��a����,��Gx)I�J0֘�XF؇}�)�� �#�],q�`_J�D�ᒼ�|���W���8��4��Y||@�m��C+�E^�6Y���p����S �"�]�Jl�0�-\�E��>�7r��<[����;9B9]��CHc�apsQ�IsS�.�&�vz���b�;��D_�Ǿt�
�ȭ��b��TG�(jt�� ��.�ϰ����/�y�+b2msQ;����v�|���>����n�Y�c{e8ͪ�g��W�~�io�%"�+4��E�r��N�+��E��? �����ijހg�Cꬨ��TY)UM��?�2h�0�n:�q��4���y�9ܘh"6
�1���d�f؞:r��~�W��ѣe�]ւI�����#���Tkܫ}�I�AX�X�!��l��r]t��6�:�r�ny���e�r�0Q� �u��c�2}�f����W�z{RF�_���+3B� �HV��L"�sZ#;�|��~���kR��W_8�pǟ���뽇���,���BG�'�!���m�L8�˛Ij�ݷ;e�$��.پ�U���m��n�*èˢy��:���y�j�;��rOL,#�������B'E�Rڦqn��%�fa�w ���'�Z\��u�0�9yUW�n�2������]��q �j�`Ec��9]�X@�`�v����2��K׮č��<����U�e/׼ʅ��D�ʮ��]�����GG�����T���ػ���s��6oMn�@�7�P�z�*����k���W�3m�.��2:�$�g�}�����~qF	e�hl��X�P���Ġ��/�s�/"���D9}�s���˕�&�Z`Ak�Nw���^��˰4�,:���eǰ��َ������[{"�f���1�Ș��햺a3\�t�e/Mϸ�{#�!�{��u�|��ĸ]��2�;�}!�i!-���n@d����S/j�(i��w+�*+�~	�t�-�i�c8'���+����z���������c1���y"��qx�cg�+�Ǐr�p9y�ly���r���-.���$���π�Wi��R�5ʗ��א
�xuӮ<����s���4�2�]6�F���R��$�ӷa[�i�}�ߦ $�q`hHYt��*^<�]�f����}�K�Ɠ4����{�9ɾ�C�+tD�ܸL���!��Nr�䅛��o��r�:�� /��'��u�E=| �Q�w�{Ͷ]J�tT"h�n?u��?_֖lb����6_Z\��`����B�����l�fN��(�Q{�!W��mv��j�6^kP-�Ɛ��.����;	ri�g~�g���
��\ElJ桪��{��-�'�)w�yʚ�j˳/�o� �i�C�<Z.s����\b_ƥk�� 4&����sM����:��n�{��D�94�����:>H3���Ç�}hk��壑ր��,��$T�����0�ց(�v%S/�J�������3L����۵n��H�Ν+k�9�|��r����CW��Y��2} ����*�!U��z"�f�9�k��j�gx��z��ba�n}��s��񡺵:��g_�=>�Pg8��̛iv�-x�����`٣���ej+4XƬ�i�q��g�D���K��+E_��̓��0�[�E� ��������̙{}8��a�����s����9��.g����Ʒ<2����(\at�gEs���@4�i)��?^�����;0`yُ�7��Ȯ�� �pc"�������8Q����U/�߀�wQ&���o��j��W��u�g1Ǐ-��=��mwvЁ��n�C?x�L�f�9&������_�^˪�����<���P7/�6����	�k�l����@K����K�C�/�7�YgU�1=�V}y����Vw�[���˰�я��S=��Ą�`T�E�N�V[Ѭ�z�Z{N=û_�m�����ۋ|�k��B�?��r(�JL�\)�}��p^��Ξ.�O�D��U�9ͫ^G�3y�$�ο��$���}�;ʑ��+H!�3!��_��+R[v2�I"L;v����L�@�`cAyy�a�^$Gb��-_���P�m�~�J+����� ��	��Tש'�����	�M�4��8�4N�:�$�-R<�E:����.�a�>{��2�47��v�X(�i�$�jl#/�m�W��6PO>T"b"t�Ni6��ڲ�����P*rL�2�&��-o��<}�/�������I�_4 �M%b�_ڳw�@�0���O���{O�<�n.f��'>Q~�d�����@~���'���5�2�:��$���,v�~�V��=�t�^z�<��K����/����x5Ŀx�f��~	���[� �N�kN�;Q����~ J�]�*�b>d��5L����PnE|�L��7|���y����ܯr�������8��nB՝*��g8�t�C�i��o}����+���o�x�5.v�_3EĶs¸C%�J��6�u��"�8�m�&��m'��/���ŗJ�K%k��R����Oݟ���k�ݢ��:��r�P�rsO�*���гb	�6��@V4��Z�T�~ƕj[q�l�=={�1�q�����s?�s��ʅ%*�66��v%�?������w�Sw��,x�/�zyd�׾x�s�G�����E�B�vʽJc�܋ �
R)��@Y�I��`�(����CDs�A)�h�R$���S�J��{Y.7h)֌#X��0��@w����O�>U��ɔCls��-�U^��'�;KY��o��|����*C��W�&��%~a+<���r��G�9�����R��z"v��AuWe����~�_?m�V։NcX;>>>Ć���>��%�N����-���pC�/OdWi	e�U&��m+��U�;�5|��� �eC��C����L�S�?��?�����}eY</�ԏ?d��Ε׽�Ay��w���@F_I�JB��g���sϓ�v9{��������;�׽]��{����S�EQb�aѱ�@.���^6�TI��I#�^q�(��:wȼ�L�k����+�n��JK��bXW'}���h��\l������,&ѹ�!A)�OX���:t*�-W�y{��#�!u��Y?�j�4���0R������Ȇc�l䷧�?�����iy�E�ݕo�l<��c���u�eЁ�̓��y*&D!]�+��,T��Y{T����'��`0�At7DR��:n-EN�"�|������h���"��eq���r9ľ���J!z˃e������/3��s��+���2U�T�r����}��W���ʣo{{��O�w��@��R9���1؇c��:݄/�ϲ�zJy���j�7+� 䅀2�X�����<E��k�O ��K$�ѩV�J!P[��r��st��3tVz�Q����tF&� ����w�� ���O>^~�;�o�+�"\��)W���8�?�d	K ��[}9[��R�9� �=��Qu��\$峝�#�A:;"����n;�p�'+ٴ!�hñ����j*�[�Ҡpg��X������ڢDuO�/�����o=��J�2�Y[Z�9񥨹(
,)Pl�F��h���滩௨�* ����Q�����n~u�M��G�/��/���/�}�S���P*�"�3�z,� ����xac����o��R��GˋO}�얃"�#�tVHf�?^o��o��x��c����O~����rm���9�0˰��{._��mNf��/p�:,0��#�N� ���}��G�ܼ����"Ew�ɖx�G�}���(���,^[���'H��R����\9���{����K/���e���f�{;�+�_��vKݸ�\{m��b�{��]}0n��K�hC;�vf�-\4S�D�r�vg`�yWܽk u��%���B6>;�~dİ�Qq�Z�D,t�ӳR��t7^�B)2�/Q�	A25�.�p�=����c*<P���"{*����}��������r���${T��:Q^ϵiKW�_|�\�t��G�Rϗ�\������w�w���l��'>R�O��2l�
TR6�rm_Cj�	�$�f"�`cr��I�`sJ��O��0 @�N��t�CƼa�MU�~��s�Pec���7�8�����<Ĩ��������T.(�c Q^"D�An�����M�m <S"�~�T��l�����ƻ��M3��5l�,�z�%G9���u���SǏ��ulǛ})eٌ'���M�m܇�|
�
d�J����nW	L���~�Q'b"N��m8������>[�����_�诔ӧN����sL�\ق�MA=�{�[�¡ٹ����!x�w�G��Λ���Ēa�:y�{I�p 驏?���>�Py�����(o�?�����3_���PP��T`���i؇MV&���
�<nݘ�S��T��&�<:6³�y/������"��\g�tw���HM�����P� �U�"I��]�  vÒ�M&Z�+���7��s��t��鮞�0���6�s�cƉ�`|l{͎V�s*��r4ٹ�{뵻N��I79V��T�$��9���;
�"���B}�5n���5NB�w�R�!]�D����r�r�k���Ǹ�b���(�Oo��G\�F�D����!��}���������,�²<r��p�T���/�0�-(���j9�}	��9&u�H������3��7<ZN������ϱ�jy�=+W9�ӑAhw.��ߌS�O|���o?�ˁk�ؓƔ!$#��a�U}��xI�����L�(3\J��u_���T�������r�����Q��2�F�щ�� J:���HD(����~4K��ٶ]�nڍc=vS��}�9��:���
G��閺��Έ�%�_���.��2�d�X�~�IFD�~E�3Q+ڧ���fX�0�����=�*�13�#1pUO����z���P�����py��'�����~w�+���,z�y˛8�vo���*�s_*'9ox���T��^{����8�����ww^,�Pko�;5�t�*'�,XO������JN�7X��D��{O��������0�T�-+�$�}y�I �`*�d.:��p�m���e	�"�����˧^:_�g�<�,��ѵu ������|�+��D{����6���7��z�>m�������eZ��eD���s1Gd�c�$}� Tfo�o�LV�P��5
cO�*.%�PVJ�Dm�v�ڣ+e�2nW"�3l~I�[~T�(�tDr�wu�ӽ���Nr��;�>����������Ky���P^a��̜bE_O@��j�Uq��c����ڲt�Ry��,י�=t��6[cϟ/���\y�����پ�P/=���R��4���S\y|����tEE�PLe����HƦa-�^8_ƨ��������#G���'^g�u�P��Ti�����,{ş��/�=�)�!۔�%N�ó���
;;��x`J��H�D)���^�j���2TƲ��m�l�L?۸�f�4g��eq<6(K&q8|� ���Z�/�]�`ȑQ�cD�cI�m��ր�6�֣Q$� H����&�:��u���K��d�!ܤ�]�'�\AK�o����_�I����� Y'@��b-i�����sr�0HW�\)/.�䩻�r���������S/���@��*w�3��W��*���xq��O=E�&Fǡ�R�m7bQ�gΔ/\潝��[�	��@�ˤc�fZ��vO�-��MF�g��������֗`n���QaE�C�GϤ��e�tY�4���(��@�m��6��-!3�n��6�Ե�M���R�IħƗ�O��xE,�\y�[��=����7]�j�dV�,��d)�L� Yqu�Cy����WU��I�w۹Z���_�i�*%0uo��-����7�jG��.��|��ϕ��?Y����P.��ܸj��+� ҆�(�E�A    IDAT���gN��P� F@����l��<_��c2:V��\9��ܸ����7�7YhD7YŜ����s�8��H��YB|2��� ��-f�7�\//r"� ��g9]j_a�:�H�J�ݶ�9P|�R�*,���9l�:�УW`a\Nw/]tw����<��LFzx�B9�v�ֶ�0�}����[���]G�8^��.��h�2o��{2�6m�p'�ԺڝTJ����ws�[Zb��fp�����_2��E�xG� YH�Be%(��-��3n�FI�2
�Y�qK�3�a3�,��v��cY��o��<�������/�{ j|D�Zd&33�/�\�>�p�v���G_W^�_^���ǹB�Jyy��ԋ/�3�ȣ0�;�\ִ�"-"������(��DP��I�D�� �_�I���/�/Ҙȴ�Y$N.��s'�[sey�4�i�ʣ+��H�ZفAp��8�wA����͆w�U�-�.u�(%<��g��C�ݯW�_�E�T5���*;�J"���aX��{�`�����g�M7��g������s�v<+�.%Me8�K��=��3��qy�hYrÒ^1��5��PG������|}�xj���π�����o�x(�]3R�&��k�ȑ/Bi�.���+�)�꯳��g�=4���|\(���BL(.�RzՆ�A�oe��!��^���N�����?˼Ef�'���jlB���N���1*娓/+�Q�jV !P�P� �Qv7-��E�t4�.r�J�vt�p�wR�ak�^!��0��p�k�'=�}#�`#��ٙ�m�����b?����8�ߎʪ �
L����H@=�e�-c�7��K����9��� �=ٖ(?Q�5�ye�����?�+�V��?������/������K������\6���Y��s+�<o}�����,�\�x��]��B؄��2\:����{����8�
]f�HVa�S>_�-�)?����,���m�.���֛[������t����%j؜����*I����aGb ��n�!aM���dK�xm���p�2��8Vw�T^=)y�9�T	�ԥⰛ���������(9X�JOr!�s�4���-�,��_��Jܪ��CU��~�'p�g�8]T�Ja5�+m8K�JQR�ǧzt�g�Q1�8���>�ܽ�o�D��f���L9�BϷ������.���P��Y�d���{v��F8�
l��8M=R&���M��a3L ��%"�w�xY��-�ܩ���9�������{�l�E�~��O�i�]��4�#�cJ���Ò~���A�@��ZVb
BB;�xȦԡ���*{m�9�5Sݴ�@n��e�������}��3����zv�dKL��wQ��w+ ,�)w�}���J���BJ�3�(��
Z�A�[�K��V�\���"@b�F)��m����O�B�\
���}cg
����=Q����o�[�ϭ��Y�[ҼMj�x^�C/��j&��\8R��)�t��N�
�TX��8���D'����8ļJ�����7�ȦsP���ǿDIή8�D<���r)?�c�Z�ۑ��wU���Oص�4�x�*�OexS�El�j�ݎ������ٸl��㹣úmno�o��*�\�)�h7t�=v��䬻�J%5�ns�ͤ������4X6x��E&I��V��oL#fU������4��*n��X^gy|�\A�6��T����_�_����?�}(gO�.�؉�؛��6�U�a�;#u\F�� "a�e��]e�F�:�ԛK-���}�r�ˀ���
K��������� ��\�:�&d�
7g��bn���;�����U��;z��E|���N�
��'�/��4S�|�Jt���闝#�m�h���N���a��/����RӖ1萦:���o�D�8��u������E���YT$Wea�2�V�K����5n���]��7��)U��6J�ku��y�SDl�1{����h���r������nб�UlJ���'ʽG�!?g��[�=�L�;o�\$qQ'������y����4���*�S��Ơ_��_-�!���>����j�0{N�fC�A*�{��U��u4�d���?����RA�A�dī����a��#ᚁ�S��_�/q�vl��]w�2������#\�C�����>�����;�(�cc��½��hA4dO����UI@O
�G�@�:dIa�~-(�w%M%�<�T���wѲ�����&�3d�6�����J��O��[����N�����_����Q��F���q��{g&Ƽo|���?����E�;�I����=�����+>>5����F�o#�dס��^���� ����nܧ�;�_B�?��ߊ��D�t6����X*k��$�҅k E��7��j%�r	��u0/̱�K��Wa^�"&u4���?D$�"�m�"y�v0�TPwyQW�iƓHU���ŭ��zf:*�o#�v�$ ��O�DV�qC` ��!��>�8�5b����6I�һDp+ 5��OVl�������a�צ��n~�L�%E�R�'��&u�Ke>;T�3�Fn㛮�<s��/������gΜ������c������Q�ao���zZH���RVH��Fc������O��'�=���(��zjh�b�5�}'4��v=�~P���K��Mi{T8d���]R5|g	���j��������5t�����@�*���c��+����ddן}#�� )���$��m��k�y������T�'�X��[ [�[�e���i���	�L߼�O�����	��O�LO]������5l׸�3��|��T���g��X�W������?����q�i9z�K{R����'��?�٧�ɞ����ܕ�G�h2^ ���Q�`�Jn��d���kOU���d���!osIus�.�6�܇���/�t3�=u�f�q�!Ѵ�Sֺ8�S��e�LYj��!�^�����&�*���^J�' 2ܠ=��&r& 2^��l����[�5~G��V6���t�e���]}�9�F����'91�UV_�����^�&⎡Z9�2+�.���쮄�e�أ�NӼ���_�AӆKs�*���K�);C�XTw�f|]`+?ߔ1è'�mz��[?�ڷj���������������A�^��_䖣�h�6hn-;��g۹^��1��Oee�Z��O]�6f�S��?���xr�m�pZ5L��R��;K5��f���i��Y}�ػB�*9����e:���	}�$F2�h�և#�L�~
�q���!�1�(��[���J�Q:�UB%��D9d�z��aj}*<�/��u�6��2톷�}�DRY��S�j}2�fU�X�/�M�q�(s��Tc�_�r�az��ɿ?��]~���]���s�9�M�mj�gC�'�M	����v�\+Ry�lӫ����/"E`���ǯ�q�b��[g�~:�Ѽ|2�2Mu&��y�u�W<�s�����mʸ
Q�i	��#�a�t��4ܮp����\��D?�������0���WOs����nβ�u��8qmC�_��nW=a��{��͍�9�jaÞa��	7�(`K����j���E�/r�k�q3��Eh�68L9���값�e�z5!0�7Ӟ�U����O��=�Jaz@H�Å�:��L+�<E��V@s*��{�{=�m^��Zw�&�K������IŅ��]%q|�����=(�E�-R� jm���f>UYa�/w�+˨�#L����s�ѱ5Ww;��ѠYN6�2~��]�4�Ѫ��`ڪ��^�L3�kX�Ϩ(f���x�bBX��|v�Z����ԭ��Y�xQoF\� �ET����Ut�rd%�?+#|����&� W�A�_�N��K7����4��^�2LX���Rtچ���a��u.�T��3~WB�c�l�k��9.I��ӓ醷�,�z�!�,z��a#r��{���i6���0�M�[�6�L�����X���c���6��v��H����8ER_݅�0�5A���i�}�P��-����Tְ�"ւd�H1�ʤ	�@�_3?=ʙq����`�K	s�gx�צ��*өY�*�%�����	kqj��%�8d㛶w�YW��uO����7i��g\���n4�x����7�y�����E��dˊĎ�Z�
�d1��e���F�rZ�N��V){M��n�~������~��!I����	��cG$�m#���,O�j��Զ��^?۳��>t�׺ny��j�������<P��\,�3X�l]Av�o������w�K����x=�U�~Z���O�aURݍ�]��W@��5�z?	hv�[;� 2���0;��������h˓ygw��l�:f���i���?��iԑS�֞�|��nYu����ؼ����9��.�;B�=��{��#w��l��A����W΢ns̤O���l��Ӏϴ� �*@������5L�͘]ڤWӼݿ��2�l���DTA�n�'�i��=���O�~�K&�R_+��ܽ�<*�J���O##_ޡF�%V�L����9a�{F;�����t�������p
��̷�g�M=�(s���i�k�$[�9�-�s���޿�G�zJ��n ��Yz_@G�q}c=��d���D6��}�>���ަ���N{�F�z��0�Gu�#O"~���Ks=����Mo0��t�fo�ʹ��z*�U�ƣQӬ��􅁝�v�~���2��oX|{m�{�G�D��2�o<�-^]D�?�q�2�w�aP�7r3pX�!2��^�
V9фb�%xxL�'��*����t��v6��&P��<X�eG����Ul�x�=��|��(�e�X��W�u���������&Ŏ0w�A�Y��0���D����L���MЮ���X�z�q��Td�)��C�H��E?tpHa�k���Q���
��$��4#��tLCjN�F��p���k�;Ŷ��#��ͱ�q��|H b�k2��_��V��-��6`g�t3\�u����,�q�Ӛ�f����f���^�$�ݦ�n;C�mm��,}�j3�f�����6m�m7;�_�׬'�:_=?�I�����^"r�g�A�iH�UN,�_]j.r��s���Sn6v��ٌ���w�I��j\wY	�Qx��-�tEI�_��T�O� p/섉����l$ː�zi��|L�0.�QO�;�2���
�n�1�{�cJ͇�u�IWU�q�� ;T�	wEf9vh,��Qw����6�y3^��()�n�XuO<ݸX8*��Ȳ���!D��-¸hf�m7�)��q�46�+���*�3�����rM�]T?ջ��(�p�9����@�֩qO�׊1EV$ۚ���n�3���~ o B�8����L��Ӟ��l�	t�U5(Z�����ʙ�fy��2�H���8�ӎ�Z��܆׼��`X�Y6�e�S$g:i�-�-4믞f���a�n��mޙ�e�J���
'D�j������M��9��[�3��K7�	(v ���r�?�S(�h`�a C�.�36��į�SUy5�J#�>u��4c�e�"��VM3�l8��'����Fna����g޵�k:�Qӣ$4��1n6�øď�&���$�
�KMK���*��y�Y.�fU_��Q4Dh�l�q�WF�яol�;]:������xN��6B����V�.�zv��I�)	2Y~��l�?���1Ľ$�1b	�V�|c»1	3���L'���>�e���;��} ��Z�X���\.ͯ<K���Ͼ���,Ö+o���ڇ7�7��F�i��=�5���V�M`�/��W@�n��+�J�0*�UO?�M�C�C��/_�?)�e�Mez7�g�,�nqu���ߦ�_�������uw
�����Ջ=馞��D���,QVt���u0��:��I�gx�2L/==Q�^�U�d���k�s���w��W�^���:@��>��������,�x>�������W��=v-�Ҝ�H$Ю��T��n�})Ag�A�#T�g7 �f��;��Yw�A$FS��=�n�W����4#�.�^"{�4�����K�g��Tփ/�a@�{�O�f���Q��mq'��5t�0ӱQٞ	�-����i�/˄~��U1�tW�I�-���ԍ���gߔ����b��Ec<��}sbj�����0�N-���q(*KwTZ t��W�h�[���Ġ����z��O�q�_?�2�l�A�tϴ�[s��b�����kˮ�/���ɊDZ����]y]hD��mm|Y�ɰ��W�.����5��a�M��+�U���8��Y�{?7�΅�?�Fn6r��l��s��f��=lx��wSY/do� ���e�l� L��f�oU�{��V����8Mok�k�8:'Rg�6O�e~鿗^�!��j��d�uJ
�S{4tJ?
����� Z��1�ƿ��G���\ȴ���0�eu�U��G[~��5�>�[{��8��Un���,����"ޕr�_3�W����'O�����������to�Ѡ�B��=+�]�� �� ��4jO��[�q2��3?�f���洧�q��;����1���#�e���龛��o�i�w��nY�����-w�@���rKLZXePØ��*a�s��3~�.˓q�˯�O'㙗��i����f�ϝ;�̾w�����	��kE��k��
|�!� w0m���+IY��-x*+$���<Zq�3^\���t3ͭj�����3��gg��������j�u��#Ы��8����֫Ъ������QM6Ds�	s���u"� �T�N��{�Y��Ȭ{�k��W�����0�����ޱ.�^��4�|jiq�WW���^����=����>=�������{��Y��da�SY��J�_�מH�9��f�V�٪������3�v��~����2L��|�<&��S�i������-|�g�A=����5*��*�}�$�L�6���Dp�2n�SOx���L;�d:�J�ZV�<���'s��WVxY�(���6�yw�x �n�0�����;l�w��D�2nV����;�H�;������Z��&+Q��i'@Ե[�l����8��k�e��lt�i6|�O�uw�A��6�f�QO�O��=�S*�Ր����+O�k�]�Z���&�֎�g{�j��$�l9U�%^��캙��l\�х�W7\�Q_�H{���	s�Y�����[�M?e��؋�'M�����&��ݕ-�7rS#A6����}��\qW;(�����l�[D��$��,�.z�1,_V8�i�_�|�_���5�[�zz����"z�g�5t?����k�w�oöf�ߦߖ!��:�~��b��2d<�7�[�M{�e8�������l�}�B�ޓN�G)�hutz�����n��ۺ�
�`[=t�3o?��s�7�ή��sQ���~Y!����$�}��[ȶ���Z.g߬�ƞ�[��Q�[,w���}�[��j�v�JiDlU�=�E�گ�T����|}����i��km���-��]�i�!U�n�|!5��ȓ<�$x��"6{7�v��*���?w�S�Q�-B{@AQ�����f�x\b���)�t�7�Flg뎱aʓ���Eks��{K��BZI�Ys[�Y��E��2N��፟ȩ�ٯ��m~�� �a3�ަ�_k�<�]=�����=��� �_�u�uk�3n�հ"o *��H���4U�f�¡��u�Z?���7h�=<����|�e�2��m?�p���f��m���2�]�}#w��:�.��Ӏg.��*���r����0{���/+�{=S\�kz-u��ߡ�ׄ�� �5�ifGJ��?�ճ�GW�S"�OC�~Y]��sF��Ou�;jOe�_��q-C���h^R��"Y�$!�w�jm�ȓcWEǀ���`��0E�!BZTR�FV�<�=ͻ�����~�nʷU�J�ئ#�����Qݻʹ��ܼ����ZX^"Sa0�M�����ّ��M���۝T�I}0��(b6�'Rd��W*Py�;���|�o�t��Ӟ髧�z�k��kn�kӕ@��#ߎ�h�3����=t�&
G���Mwqƻ�Q[����q�K\I?uݼP%��Yx�:̼ⱉ��5�q��-����w�����=�ek�{}��5�E�+�K�LQBB'��T�b��    IDAT��W��)J�t��a��=���6?X	�^>]<ä��&��_��i�#��8�9/�7L�aڸ�1g�g��UڝhQ�0;x��7���a�b��q���e�v��j~�
)�69�ۺf9uKs�5J�u�C���ԭ��7�*5�=�@r_���<Y����� 2��O~�|�����!d�M.����u�;���� AQ;z`e����ʳL.��ig>�i�u�<3�z���n�{�=U��v�6��}?��13�uK�L��$�fy�rf�W����</�n�ӭ+,�=�=�gҬ����n�+��B�@m�V�i�I�7[�\;Zys-�t�FW�3�L�يe��̳"��=mȦ�w�� ��d�=��2�LW�H�yj�<#\�-�,���E�T7b��bχt��#巜���s��o8cd����Ġ�,��R��*#:�mq߉&K�Of�6��^8�~�Qe��}h��ݩ �#_k{�L!��ʔ�)e��ŝ�H�E�M;^G���ޱn�*�h��Ӱ�	��?w����V�G��g�c<���EI\b4:��L�K8R��g��ݥnsParb�[1��Z�������A$��U{ �^��'�5�t�-���8*��LO��m�̣�����3�;�J����S�3H�߽}�3M�����Z�#,���_s�1ӌ<��+P�z�I�H���!<1X��b�~v��|��-ի���9�n��;������1J�����Nv϶�fE+8'�@EW��uo�����=U�����=-wԓ���Y����y�n6��=���[�ߍL4�v�z�g����n�NSߌ�.��&G:�~��~�m:m��%�h���sϸ������[�iʘ����I8݈w�m*����L/�;�u��}gg.&�y�6���[��u��-c�ݔ�6�)d�Փ�nF]e�l�Aզi�L#�����<N{���n��,�ni[�TmY�m�8�e��O=㥮{~�z��7˒a���ކ�p����n���f�Գùx�{�B<�kO�K+�vK�u�7�f�,���
-�@^Y�M��`Da�{3�Gg��ߠ�J��e:��ֆ��9Û^旺n��n�{k6ܗ������gڷw���zp��x�յ@��n���.p6zv+�vsҚDG�b\�F�^ڤ��qSE=;Xf����'��Ӎ���CA��e�fK��KoY������U�������p{�w8��E܆���`��˟�r�z�M�
��n�m�*���	����i����2�Aw�;���պe�>�_L^6�z��i�g��~�M�dz�iΰ�[��F�z.��z��{�sl��(
\�ۋ/"�^�b�G=��G���l�ѣ �C<:*��3|l�,��\�"�*$��z�`�X���7��x�q���5L�֚�8m�m�/�l'6��2=���񮤢�u�ޖ+�Gܻ�؆������-�H�{�5�6ˮ�O�yd��=�Ͱ�u3|ύb�(�̸���'N�oO"\���I\q������:�k8��/���,������
���a'$^Gfa��<Se�'`�-èO�a4���n�t�4RL?�gx�v�F�KUm��&-�[�^�;�i�i��:�W�5�o/m<��0J�D����<������"ͮ���[�#���q�r4�a�<nܨ+��}�˼�y��>=��=<���-�l��. �������1��mʱ��@j�WP���w�~-r�/+��L�Y�4'�ɰ��f�m�~m���p��J{�մ�qSe>��Ꙗ�6�iti��ƕ27YGr�g���tul�O��[����]{}��Բꖓ��]���~v�]?���&i��7y�t��m��w.aڙ���'�3�n�;�����
��#�w�l���g�l	p��J]��zAO��f�� Q��ůV�/U�-�f�VY�T�P�3|����7�N�_�q5g|��9�͸�e�2��K�0�t7M��k�2\�����`m�����o�hnå�n'��kuˬ�1^��a#�9����X>�M��/n���=.6�"�8z(Q"'�۩,��9sWܽk��2׍L��e�d�FdFq��fȹ-[�z���]�X�p�,��Qw�*�����ӿ#i�m���2�id�hT�����|0f�W�Q�Y�^i�ѽ'�Q��t�e�p�QJ?�CM%�u��xY�t�Mw[���W:�|5e��{���OЌ�z��G��=ӳ�!m�k������"t}[�����k�q�[fW�C�܎E>�ޟ��*��Nպ�Ӭ_��ά_����=��O�i�kW�g�p�~�=�w)�H��R��}��F�rd�3��gg���ʶ#���D�����L�g2�G��+4�����0k<���ӽ ���O���D9��rAG�ۓ8�F��~w��M�y�A����K��6��Q��݁�V`d%�0VZ5<��g�3G{-�&u�MՆ�M{���n~�iؓ�*�ɖ3�o���~F�>�^c�{��i��M�L����'z������4Y�V7���Q���42^��h�n�4z�3���Twۢ�����ק�y1-ٓ���a^;H�f����FnX� �vS�h��?�k�kX�Y ��~[)����m��j����id2�`z��N�_v�to�[��t�\9,��_��q�4�U���j�Y��ph�N�֭5g�t2�z�k"��;�x?�3G"^�P�|ϴ񏉦q�s�fN$��m�m쒾��o���2 �L��`S�*�ʡX�D���pP�D{��=�5n��j7��~�3�t�3�tO��z�%�ʔz��x�z/�@����3�i�{��@:�q�+�n��-�3ʹ�H�[�4�f���fôj0\����a��+-a��%�HBҦ=�;�����b�T����\RY7�D��������������uvj�r�����:{Q"wL$1Ǎ��f��J�f�iO�hn��9������z�@&ͦ�*�2^��a�r2�f��z���ץ�i[�Vq��gm�i�����2�F�c��/�Id8�/�Ro��*����ZQ�t�,G�A��a�H�t���(o'H�?�TE���p}M��Uԉ�׷���?�FnVע��1[��f_�D��l%��d�2��,��7��Jd�Z�K���6�u�������܌�j�~9F�� \�z�x���ȇ��꣓����i�X�t�Uδ���a�׏��{2?�T��nm�Z����F��bF<��Ong^'�+oRw����6�ʜ={o���	&FK����Y
V��ʒǧ&gx�Έ���1*a���2`vTwx�A}-���2?�TO��t�J��H��3���;Xh8��f@��Xh�$��<��Ꞅ�x�c����:g�U:[U��^���"m��(ʟ{҇�q�$i�ӮDV��7yP�Gj�sNhp��/ab�=&���IbO�o�n��gE���ߠ��>��-_z Be���򧍓���=�$d(5�H�ig&�˸�Ty9�f����9_QN��k �P��3(�\[Y.ss3e��R��ˋ��G�����́�X.^'��|˷�?�_���
B{�(8>�$�ն������/���g��BL����"��yx@�R�N�\MI��܊"�e�N�^�.�:RĦ�zv$�]런�#��.�U-�zp��R��_;��٪^x5�w����Ӊ0]�v���#�|)r5�l���8}�5\~g"�b����G+
eST�'�VWI�SUJC�p�@
���HD* )�x� ���� vT������c��'�b�d�
o�;J������Җ�$�v��\��y�^N�{��ݟ��r����Ʒ���Z�g���ۙ��賵�X�\}��M��H[�?C������~�7���;��<��3��C���%�����"8��6"Ј��DT@���P��H�b����L��4-B;B�
�Jd.��G���X��[=��ꔐ��#3�4(�%(��a�_J[A\̹�p=FDPj����H���r}/EXB]6��xfud��E�j��G�x�2UT��X�A��7��n6z�3N{�~f����޵1���W�W�B{�ڣN33�m�J98;Wn޸�9U�\^ �7���گ.����<��7��Rϡ½-Q�'?��e� �mh�^�+C������,��
^���[������ce�ȁ�|���?���W�cÕ�1oG�d�qU��傲p������:�fWg�1�޵%�G� }�g��lͫg¹�h�F7L�ӯ��!�~]v�e��#ZO5�^��S���w_�ϫ()9v�X���ꐭ����`�7r��e�Ҏ���C��#��7͂����S@:+�[y�k+�@ɰi���q�EH�D��=M^C-�ٱ7��9�������R�n)0/_�P&aU�a�W�ڟ/G�,���@�Q(�X����z�*� \-˜�C�A���g׸`���h��5̲7 �ƭ����{�3��w������r��8��d�yG�/�o�*e9G@~_;Du ����o��� {e�R�@�h&�����'�G�5���7m�O�F���_m�l�q�)�!��1���F��N��B�l��������\�w'}_����������$������G�`$�L�F�2���-��#���h�
0+�{ �:� �v�!|�����>׹���ި�5�y���s�9��Ux���J�k�W
Ѓ績k�|�w��������׃��v�
H3�q�	�h9r��L"���%�����8_&� 7�Q�����́p�E?u�^�|
~��B���J6�*����4�NԵ�@�pՁs,���z
gU�b���֝�f݅M��]2�����_d�D���i��e��-ä.��ٷ�5���_~�r��щC�N�6+���=:>�q=��9�l��y#ޥ��y��Y���n�VJ-"��2\�����}*�q�*�@�|)�ʗnu�[D�0ye��0It�͛ 0�~�W~e����r�� �+\�?_�^�ä�~yy�LN�����ū���	�ݙ�aX�_�l��
H�y�3X�i؏�7.�q���^)K7��[<lt��da?|����{cR\�+���X),�p����p�}�jV���]������Cs�^=үI�~��ԺB��Ʃ�4�Î�e4�NI8Uۖ�v �;q�D��U�2�i��H�2� �wQ���/���wY��q���o@�W��V-)��[� DB�.�Jo)PV�F��dD�g8�2l�Y"�@k�䷕��_K�"��[����_*����ჇA��r`�`y�����q�M.i��ˡ�sP��6�a�౫:�/߲�K$¼��Z��)K�܌nL0�X}���t��\�l��ó����ꤏ�����e�NW[�"P Q :YH�QN��ȦN�D��	�M�
�|;'U�*탰�=ag��+͉�3R�'�[�^(Kg0_��{��c�VWE�*�
mż|�Z�����ͯ�X�����7֜Q�ܾ�><�-�D �t\j��������k�ʉl�J����D����#eowUk��,���QB�%[Q��>6֟������[ʛ����	w!�'U�2�E���;EF%¾, ��ZE��X�>�V�ɩq�?T���4(�fsk	^���n0�^.�`T���T���(������J�VaM��� G�B���+eb��:���L��ӫ�k�^�� `����#�^�nP�32`�|y����R�P�	�w�{;n�)�1jG�B�)Ͱ��+ݮ�M�]dh�ɱ؆B۫-��rk���~�j���'w���}/�/�]ʷ�l���^�5�j"����* ���q�̊Z)�KU&��>��Ͱ��d�Z��5|� ����N�$�ȑ#�sD	9�,�d,��������<W����,��+י��bbe�7���2A�SIDuK�e>zll�k X����v/��$�-�X:̱=<�F<�G>;�oxd�,�|���C����W*7�/��).��^�%�����Ab�$�� �R�	���K�΅�=��������O�M�����m�,��(}�x	�l?��	�#/�vݢ�;��a"@'����o�Éz� 6�nӔ����	=���Lp}_�}������u�n3���8�r+G����iq��ʷe�0�%b'�w�%�N��_��]�"�i~)��q�A)ȱcG�&qR����K��`�u_����Ώ� �*��X*d�1���< ��fw�1�ff�=�,�CJ7_+�P���_����cz�S%���\ER�� K���,��vbb::���f��*z��Dy��3���.��(߶����Vοr��Xܠ� -�.���9ne�E��x �λBgr@I>��6G)�U�_��#�}5ؑJ�T?�;��4���ILG��໵�YK�	�1T��<R�9Gn���m�.��U>��v���ܣ�ܨ�bi�.-l�,��������e�,`���+ ��'�&�G�L =�t��;�2h����b���PaYCj�p��bʷ}۷����{���O���z�I�*7v�ƅ� �K�  �敠֛KP�eq�2io�C#1Y�	o�L\����,ȸ84�����3����k��.W�!����]"��x��2[<^>���r�)�p�K�{(�ty��O�����Ay�%��	D�W��,Ӂ&�8Kt4���I��� K�D6F�4����p�3L~&(r�%�U6ݴ�T�q���Q�j�I�쬟��B9s�yF�ҥ�V�B�6�%���T�zcD���~7�xR����;����5��m����Hs���ƌx�V��~����0�����wѝ����}wy����C�'�]���ϰ�a�.�27;Ų;T1����-X	d��S��˅K@d�h�B�^,�K���k��LM��	5�Z9vN�'�2Y����30cS���	�1�
�W
���������˗��O-�_\�,o|���#?�����?\~闞$}�X;������M�׿��
�p�e��]�1��ا�����=H��P����v�&��4�t����6��{/��jbb$ؓ�����c�������;��ω�R����5�غo᰿�E��Z�� �պ��
��h��WO������ęu�y�zH8(+���޾���|���E�9� �6����|q�I��R�m&��K��U�����}��O,�l<�LM�Drb	ȑqyB��$4
��Mf���,)S��U`���H9��e�ztd�:2�y�tf���rz{�{˵��'˥k����ϗ�O�����~�)��{ϗ��?_�|��r��[�|>d�#�[g ԃ�bP�@�mR���RdV	����?�t�v��to�N�ȡ'çn���/:�fG`�\�9~��Ёٙ�龗ڽK����"���6��GJ��F�xR-�8+�%
��v�|\_�d�������^�5�F~�b�.J�=��"�
��р��n!~��^`�������o��߈�׮]e�u%�k]A\a�bhg'��B��SS6�|y��ϗ����@��P�u���ˡ[�c�����/�O��2;��n���V��C��3� �#�����K�0l�ְ��B����ÓX��?�X.^�h�F^�j9��d���PN�:Px�x���|-���)��jm��I^o���<�TVJˊ�C.�+��K8���O�JJ�07��F�N��btP�^۴v��sd{ն��:e9��ٮ.�u�p۫�o}+,���q������=]jw��Ŗ�]��9�$�r��=%��\[c���*H� !nx�^�V�Ъ�c{fcO~2��4�:H6��-[��tӬLԕ�{�9�$�����������A�X��K��^�>Ϟ��@�nݼP.n�օ��z�A<�ݤ?��>�b���mxk�q.E�j*C�Bg��iD
���Q�Q��%�5�F�xG�D��sK!�^����F <bL'�k[A��M�-�_x��tu�����v�E��嫿�]�G~������b���v(��P16H$L�������4'��`<����@���v5|�W�$�팧ҽ3�8��O���1��/����O?�4���&DV-.$l�    IDAT7�Qw��Bn��!����6�׷��s{)��8����%� ����Nܤ]#s^I��w� +@ԿҲD��<��I6yE��[dB#*�0������|�W�BT�P��Ef�B^�$�}쭏��}�/S�C��rm�O�[\�R�ͯm\�dM`?��k�W���4���H����Z k��3T�m��^+�ť 9�_�ޡ�%S��L[�md��/ D�Ed���|��	��&c~����jϢ�y�b�
s�f�<�j��_|��9�@y��)/�|�|�w~My����G>�I�����h��r�nHV��I�Wa���"Q$�� �A��h�!��/ʁ���eG��l����0�v�hGe�T5C �-L�9U	L,L5!� ��Y�gy�u�,o`!i�w0�{����)�V)����{����x߀2�Z�Ae�+@�Lu3�a��HѦ��җ���"�R����d	��;����W�ǿ\���7�^���<�����Di��IDv�`]���\������TtrJ�(֣��O��D�I\�2�j)�TR�ӱ���p:�Fa��E� �,;WC�`ǕOg�`�Ō��4�PpxP|@=Ţ��`��W~�V=	>5�uc婧?K�b��C��B����=R~�_�kF�U:�WaGY�B��(����Ŭ�*�M��������n����Źb{�v�i�������ؐ�z�¤Y='���#���xrr����ȹ����l�r�=��мڕ~ƦG��:$g��Z�@�[��_tW�p��pȬ���6�65�(���I>�}�(��Y���������+ސ����(tc�=�P�!�|�������XLaG�6K��K���@Mi�\����mv����bI�JLR4�Qc�� �e��ENp�ӄi��CL0ch��[��~@�qS�����(�<����a�S<��j��	�㾧<��2��������b�|�����n��-,��Ú��P�#���[��&�3$n�iɭ94�խ�TY,���Tݶ�.Zk�^�t	q���[�u�vM�	Oɢ!��ms˦���go�/����B3~J���ۊ�ږr+��u �9U�ڳ����Tm���N 0� �z�F�ڊ���1{�,�C�>���'�xQH͖It��H9�#�^�Zo,/]`���<?0 �+�L#�'�v���7��3�dug���iT�,ӆ�8��Hi��r{�4�> 9�:t��A��!6������ �=Ӭr��3�З����3��3���}��{���CgCl69����+�����}nn��c2d�9��v@$O
CD.1��N�8�Dp�+��K���l�A����3�4�ܵ�\���M�Cح��.j_�m�ԁ&�˭�e�-����.��Bν�[������+�� ��B�X5h�תL'(�'�M�ೕ�L��</��	�x���]����!b�q�z�7aC�K+,��h�[�_)����ي���r-�C(#�U��.���1��T4� �e	��[Az(R�.����\�R]`E�.��4H��q�E7y�j�+��A��l�f;�Y�|�ۊ��cL�op>�$�>T�y�Y��\�?���ןe$�����|�ϰ�q����Cl����Z+���V-azM5ipy�:_�A�{R�����5>�̿l�a�)�S��N�$_dv$"��!N�C�&�Vc�s����c��L�븳���履�[��kkt*�?P�A��Y��l�Y�;�m���G
�)�×�u��={_9{�Y��c���D}���[�!�[������^ ٖ
s�r�� �Jt��a^�`�]�`�%V���n�YCN�T
�������]��9(�Q�8yb�r��lh� ����q���g]�f�<�@��Nv�z�_D�93�\v�i�V�)�jy�u���˧>����������{��]��O�83ð)�#�&:L�6	�
�7H�c1P��S�Vm��aj�D�Ԡ=�S��6V��e9c��+��`rw}_�mRtFI�⿡���IVo�T�� k����*K���	���H��2�n��6%����
�c� ��~�`�{������C_em���|���ɣ����x����]-Ǐ��� �A^�^Y�H�r<�emyj�r_�����&���A�`��g��J#�&��Ll�E�>?|�<�0����l�9��d&a��H+�;��/U��}Q�1)�n����r�=����R�EʽȹN�K�^~�W~�E��r�����g�/�FD�u��1��G
U�O	��	e�~�)�A�У�$���� ~v��U5��K�V;9 [��&�@I`�V�bK6f��N2A�z0��j�����2T�;�(Ȗ��ٹ�J��Wi�a/e�2n@7�v�A�o^{7�n���m��w��]��q���ny��s�M��͛��~]d���ؔ�ؓ�����Ԙ}%"�Ag����xk��D�Q/��	����@��5 - "�<�,!�'�0;O�2�2���Wʺ���A�Aٙ��\��b��F�D�׺���;�?�����'O���y�N�	������g��\���O�/{�1ح�����l������BS�6"J�P�%��0���ٹ�[\/���h�ʥ_�U��/�Q����OGm�%y?�q=���V`wvNLL���
��j?�=�6��6>��uxt�R�b�ZY�1�L�����iΊJ�����_]d ���gxӏs�l��a���a�+��?��7�7�K�.���W��D3l�f+L��6�巼|��K[�� 0+�na-HP�An��A
��v˪�j��ǐT�pCl��)����J�n˜f�7G�9D}-����H��������zZv�1S�*�X�5c.�PQ�/<:ʊ&,#�>�F�*��:
W)'˛�t�|^�{U�?��)���}����);{�)���F��8Ƥ��������d8yn�t�m���*[8&ǘlW)m���VEےL?�>q�6O3�ڎ��z#����ro�d�2!H�7�˽>19�@��[2BK�l �Df+����T@�tϲ�=�t��i� 5�圣���ه�._�o��U'�L8���q�E�tj�ʱ�ocY�ɛ[W9�H'�7P��e��|TJ-eID�M('����[ 7�?1q�L�jx��Q����9���|�uB�Ȧ���4��h'"q�l���G�iE���0�\2��Od�����l���&�+�`���3�:u� ��O���K�g˻������?^>��%��
�?�.���#�u"������L۔Q�"H��"L��8�X�g�<�;d'�h��,!���숬�5��?]�1+���Ʃ�W�F�U�U�c�[_[�➍z�����È���,�3s C��9j���z��k/'�256?��ᡃ�����?��������Œ�R MI���H��1�ZE|6��P�FL��s����2�]O�ț���~%�0%��h :.,�v�!�&�P�9���a�Ρ����|�o\"�u�27�-r��$�I��ᝡہ\�h�\	�"� 4�p�rJ夤"�R!E��`;:���Y����p�C�3�����#�R������Hy��G����-��g˯���('��|� �#�#�l�+�9w�lO���C��\�T���Iwu�@"������ҏ��Re���4�𖧆�hB��Ǧ�/��?���e��*e�d�}��%Ûc�l]\ZdQgh��tH-X4J�:[ɬx">5��GEDvT�	�~�|4�p�p� �,�z�;��w�}����G�S,\�����?8;�􁳍����!6(�k�8R�^������HVDn��lَ*�ˋo������,[��{7�/�l~��+PQO�ߢqq�L�4��9 �@9��v)�&���v�<e	lt	��nd�"�Hb'=��D�ƗU[^�IǞ���eo���R9{��r���m_>\>����t\&ǫ�����_G:$$�rұ,�Lě��S"o����v�uwس9EX)w}"����ϭ���2�(��Gۻiz\�y��7��^f�X\��� o ʑLɟT�r�����Rɯ�H*U�X��J$�J%)W�"�P�%�e�%SV��bDi;I(�@"@ �%,vg/��s��f�<���}=�~3+���y�~߾��ӧO�>�M��^/�v�l�;����N�ug�;.�C�=�<rnfn
V���2�`>,+oq|���o�S��is Lt ����fD��}za!V�V�n6O�	��Y����[�h#�&�y�[�]��<�6C�G) P��w�GG<�*2�=��x���恊Р�O�@�r"�}LdQQu���@(�@�J����[h 2A�Go��6(T$�8Ÿ��9׮�-��!��<��F֜��*r���Pa��%��ҽ2tO�t�?`	R���5(<�O�m��������	;�|��OQ�s��=Ӽ���L!�调�0l�_;�4�N�{9eU6�N�&�r��A�Ei�il۳t����=	�,�����ᅭ��y�fL*��g�[7�&�ve(�>r7�m����oݞ��_�=y��=o@�1H9kﻣ"�X{ؓZ���Q��}2�^��ȓ��F�?��⥋ͯ����7�-���D�}%�����NN�Dd�-a��6,ɶ,|�{Qw=�z(�,�|-lX���EU($ϼ���-��[��a�#���\4�����8���
����.�Pw��N�ha��Q��6�ґ}:��OE��҈�R��J�Ο?����u&��P�]nn߼QXf�r�?����^C��B��<�#TN$�X��uځl�X��Du�~�v~k#�滶�8n�H�L'ڟ�E�dh�IVlmK;��R�c3�<G�c!�����ѱ���	xl7q�"(�h�v
$���D�9���`�2L0� N�6�x6�1����ͩ3�l���|�cO7�}�2�bV�6���{�E}�j��M(8�W��(��E�Z^{���Ԏ��!���@�eA��	�ڃ@�!\�)�r9�t�?'�P�-v��A��;�Zw�GAN�[	�7uDh*��@��HKG�C�$�K�и���<���vXҢ�v�P�%ٛ1�?yd�fd١,7o�`)�BP�˗?м��nsE�S�G�� ]�����Oތ �UF���Wʺb���SW�;���*oψU�r��,:(u��P�@X����~�X���";la(��#ͱ�����橱����m<������v-"V�X�w�8)p �J� �t	�� �~��,t�8����왳h�-�󆼝�a�r�Qf�U�����/��x��2������Y\hΜ>	�w�!_k�o.d�SdJ��)�cL��/�%#��l��~���8�A)��.��qO�����K�]�Q��r�4)
�v4��è�dމ�������K�c�騒���,�ad��],�.4o��Լ��+4��|ꙟ@\�d����`�9�C�k�N��v�T�إp��X?M�����^��s{�eJ��[8��H\�3���<Ta��{RW����0�Bp�]Wwzjj�=��r{�ܹS�� r�bpϸ.�R8�,���r�n��}מ��]�H��t[ʪ�H-��N[����� �V!�qa+XB���H��,γ�`��.��;�B	I^]Ʉ�>�urj�F8�t6�~��`�%��f����; �c��P�R'T\���F79�O��&�j ���K��t��u�CV����+O����� �n�����:���������&@��S�2k��.�9����=�D��}��?��\�4È�X��g�h���w`=v��'O7�,,�09��pb@�\��{ �m�[>M�A!FR|�=Qd(�3�H�J����㢻�p�3&���i(�v�8u�D�ХL�K���s+.X�#��� � s,�F]��eK0F8Df����3g�R��8[�اPD7VD���"V,�
�����6�t�h���z ���~�s���.E e�#�@�[��i"� *�Y �P%�(ťLPKQF���(ϩtF^��E���s�߆�B��6*S��vq�C)Ï��l�*utW��9�;�T� :�?� ���v"(7��23
8y �B4��x�?i���n��eP"۲ƙ*� ?����ls�6#�D��gcʹU
1���5�T����=��o�y�Hem���2;'��3�5Ri;��̢���s���T��⋝Ev��#��t�g��Q5:Jav�)>α��H2�,#��q!5�EX+��n.jԀ���E�|7��J��|+�8щa�s��_�p���[��� ����w�fc�V�`I�*�i����9���4>��{�ܹ�w��|b|�Oā�kk���e�1#���AY)����Dh��"�R�Clޣ��bv��<�vG�<�n�ߋ�Zg���OJ	B0B!���F�d��S$'t
�-�-/��Ɏx�2�_��:2�A��ANB-���6�Bn�����D\��2�n����.�?��E�9@l�[7��G��$x��ӟ�bt����DsJ�����@@�h�� âǖM�D�a�>(C�=R�3bL�����6 �N� ��&=M�~7��{��C�C�2^�� ���ab��U��,�#�6�?3�s׍TT���A�">*�p	�G������˾� *,M1�3��B�-�JKm�jzuR�P)4y���a�SyT����OY��Ő&~�0mt�B-V+	�>��&:s�@�6v�F[��03�����2Ɗ�"G1{.�;�pz���a����˨K;ʘ�dގn����h�Kw�i���u1}�vd�7p�#v@�}�+I�m�ӧXu�И�ixD6��:�.t�+]��Q<"���6(n�"������X +��P��6��ɰ��nCGÙfĜA}�s��|��*��y;,r�*ɀ=��4�i��md��6�G��eؖ�s�
�����	��ὧ�NCV�:�/*$M�3]<�`X�`�����*�pQ,[��ٜ�Dը�ҋ����T�z�伌1Z���Pa�O�Ex~�:A˦�iB��N�B���O]H����	��zz�6_�o8�������Ia���Ňn�����z�6eW��ZPT�m�)
ʻe��R$�)a�5~lߚI�m8�}l/������(Εr{�T��4��A=����@ü���,3�2�x������z�-U#�h�~����)ݲ���t3��O���5?��?��;ɋ�L��Q{��Zmבּw=&R�`qup�����BcE�@n5����O���a9"ɶTY��O~ԣ��aQT��p����ގIY��A	��^� �E|'� �!���E�^PVQ>\ � �[�-�CG�I)��0��>�(JWv\�"�^;�����7�L�u�F|��ð%�1t;�&a#,��'
T�DhB�����[�M\H�D|�h��=�Ay�˗/3�,2��'�Rn���Ly�١8|,ʽ�>�a�/z.Ƚ��||{k�}���VB"t��pZ�Z�M��=�Ha	��1��=�я6���3���po����!��q�0�Yą[��LaK@n�;(x�0�LT�%���F��&��p���d�jN�jr�4$����u�=�L5���!m��=ؔ�oa�L���f�!l{b�8N�4�$���AVo<i�g*O�\�4"�=Ԓ%7O{����T�=�y��ع8{�Dsay���'�bQ�*�֐�й��`�P-���c.Qnʐ&�F�5�1N�ܸ%���p���Ύ��,��jwr�B�*���kK%#��?�b�����ʕG׸:a�.JJ ��ʘ���!�d}a�7+X��˂g�� �vI��[��E?���Φ��=�� Ԁv�O�=F�@L�V�3��'���|�q�ײ&n����h�}A�2��RM�_(f���ڥN"l��#xr���8%2X�B��g.�qi�z�8*��:���u/�mGa~����>ق��#!'VT��7���    IDAT9x���K������M1�I�-ymD��n�Kh�(5uOc[�ư��2���m� �ߺ�"̌��ȗ�x�)��I�]�4�ys���y_���X���o�fj�H��:�a�S��<U�J��B5��wZ��~�kچ�=�����&z�N�
�����;6J ]�ۨ�2�;�t��L�c��<�F[R
 ]��e2ʉ�q�$C ��;\T�E���M'��|�GD��	�=�b:r�m(,��e]��',
rZou��� I�~G�5��Ae<�O.,�)����Uiy�g�i�M�!���z����x^�t�#���QYF��KY�;eK�l#˒����1�������^�o�gZ޶��Y7ꃈ�+�D��0r_C����'-�3[�Sc-g��mc��V+���~[�4~�O�k..�=�I�0��;4���[���"�ڠLJ2Ȟƴ��\[�6Y�ʨ{Z�}�+�U�rƱg����l��.��ij��p��#�?���~[?��~<��'UV]�j�PR4a��8�#��^`���I+�tT#M[Xy��>R�M����L,�)�?
ז'��:d���:�n���5��ER��M����zDgD&�l��<�k	�����<�<{�9�=3) �#3���,C(�`ȑ��VW�B;�/��O�uO�����/C|� ��p|psn�c���m�ڣ,�xb��r'R��,b��%U��5:�*&��o&�ml���{f*�r�ȼBtt�Q{�eѨ+eS��kaUJ}�uһԡ�V��
��>11�[W�(����&y2�
�7�q�t� xAf�&�]�,��}<�@��}v� f�]:3������Y������v;���y}s�;2]�үg��L�{�m�4ٞ��������P������N
�������H��:���%ix�,GЍ�G��4�Bn�t�愸=A@�Y!&/#]�
�,t��<U]�Ұ}D��LKMy�%D� A�)�`'��"r����P蕣4'gV����PrM�#�m$J&F�S��S,��̜�@˳(d-�S�kL:�,�;��G�2�B�H�%{ߖ��c;|�V�b��u�*�)	釭\^�{S'�Kǌ�pTsN�,�|P7�dY�6ʄR��T�<\CSD�mh�&u���< �|9�`ƝF��sQ�(T��z��z����dq�T��{n�.�D���rQnY.�ua�j���Q��#|-�I<��H!�g�Q�oJ��Wu��"�aE�%\+������sS������N���9�do��̈�R�N����V���!�4�+����)ZS�E��{O�����sT���_RBJP!�g墦C��v�����Ѣ�Q~$�PxE}�ϲ���;�<�Bю+s ���X���u���:$(G �Ҵ�@9�{HQ<L�%��1�D�w���	�|M��`"����@�"�rq^��e"��\���$"7Α���)���Xp�����QӨ�$05�ƚ���1���n%���~�"��iҶ�GX;���+�&��:k��Y?�%8"��*{Gy�6��^h6��]���O?=�ۯ���"�˟c!7WS�[2�}@���B�Jz�����i���-i�pk�@Y�LC�E�mz��9�m�p�#�;��3�2��aC^JN��#P����q�O��T�CJ��#� E�!�pw̔��"|�˚+E���Do󑅂eb�9MS��Š���14+�Sƾɉ��}�Z���a�-,*�R4�I~����P�KU�ԓQ�i��M8����|�Evق�U�H!���u5Cm����u+�y�W��(VJ?렟�6C�u7_�P�S`/2�	,��p�V�&*����oR����c!��佽3#s���Cd�H=)�����J�
�h�\|S��~�dX�h���ïMC�ՑHJ�[��I�����I!������*D�[�5�Q�g���[���>X��j:Ƭx���N�R��AS��o�u�����<�X�$�
,��P[Xm��.ۤ�C���=�x��
e�y���oE��Q*4+��z�����d�E(�4��U���İ�;I�����5$����k���MA�lӴ-�5��&�ֈ�Y6���
R��Z��6�z��s��!�
�;���f�>�÷�s,���Do�L)��܍��؈�3�JX1��0"��T*Qz�ˊf"�?M���$҄�m'b�p .�M&9�� P:w���X�	���
��~��D9�wNs�5Rs1�o���A�b�#�Px��{�_�?�%�6�L=��0ދfb���@H �H(�k<��� �;�И�2�r˺�aw�G�A�=�mD����g�=T�\��6�E.=���9�����l��fd픰d{i�)e��,�Ɖ�m/K"�Ѷ�0�/�/�Rw�g�0v<Ag��T�Q��{,�f�&fBU�C�������
[	�O��)�e�Yx���T�r�Y�"��fG |l�U�IF<�W�Q�/�����n��%��G�����>�;\h6o��ȵ�k�p�8�r������ԍ(��.T���^���ə�� ��l�l�=���-T_�,�tz��-=��хf����oI0�Y��E�ogvW;��ߜ�*�����68b:�s��&�ٯ�$���ɤR�Pz�Z�B�K�R��%�b"W�sK���l����7�.=r�(���"G����'Ȳ��v�A'���qwCQp� �Ny
���*�j�0�M�$<i�e�
���ò��o\%:��fݼpu};���3l=��'&f����[PL7��ds�C�~m�ե'��%�E��D��͆�,��] "P�l�b���qb����!l=	m�DD�:y�q6N�h�}�D�g�! ��t$@��b�v����<���GSD�w�#E٥��;�_�Z�؞L$��Id"�cg.X�1�(iy��:Y�tYv�DjY3B��<��wZ��'({8!3�[��H"��д���I'�(ID"�".�M���Em6�N�C�L��<M�a��,]y�E���tg����y}��Lr���&���E�BCxΨ}��X�mt��1i� Z\�����t�̙�K;��
P���2i�Dj�}Ԃ��	���`�]z�] �%��J��;1�q2�xC'�HFܛ(�(��e�<�[�3��w�|�!~�C�~:����O>�6��)��:�����!F�¦�.�
���"uA�9ڕ���Pg&�¬lE#qD��ә��\qRr��M�6����n-sG�s���s�����!?�B'$��0ѹ��"�,�ڞ�!��w��v���Q]	�#k��p-���k�k�vT;��Ȭ��[>��A4��{nl����׮\9�KA)5�B��ݭB"H�L	�����*�NlV��J�F�C���\R�(	?�����6���'��&�����
��^��<����g���yW�|��)��b��=�.�Ih3�����'mHW#�����b���3��ӡF<�RD��66�&(��'�D"~����וp�1���_9�av�֊F%M����G:R��d7�,����D#�(����i�u#%+JF�7g���tf��r�����Й���Ǣɏ޾��j�><�����b?�bY!�
g˒K�h+l�Dl��aie��ݶ��/r�#�������Q���eHdag���\��^j�OI���$�)YT �'��0�FK0�N!��"k~'⚉q}�$B���;�H/��˯��j�/|!�^�f2�Ss��z""�G�y��8�Ȩ�7���킐� �M�]���?�J��m�8��|�=�l^ �=p��86�Q�] +{IP9;��@O�-���䫿���HPxu��=PQ;��шJ.����5���t|�BD���tӌ̬c���G�	������$+bF�Ng++�a�pB�-[����ͼl�|t��iDn�4��[��,v.���(�q� �u�uaA��Cͱ(���l��V�B��,X*�y������N����H~[�D�H��"�)v���{F��k�Qh�YF9��s�8qT"�D��=���8S���)�G-Ȣ8y��/�{��.G>lnrq*[���\�.��c��J��a�INS�2q��TaH��,)�E=[���i@�bS^Ev¬P5�o%�iڐ"�1�4X�@���Q��d��zj�x���v:�2�Sd��F�&{�|9����qD�)�Sq XM9J�E2�v��ߦ+����iٹ,����� X�#�1�i�蚨#�n���`A�O�ώ}�k_�~����/�؈��9r �m34	4y��:����з-���!�F��H�F	�,���G?�߇Ø�@��.qè�\E��F��C�ú�����`�;��!;���skو�H���TEv����Z�6�o"i���5q��Uz{49�-.�4�(Ԛ�hv.Y�,AnǆB�ccBԫ��2��ǑN�y�ƵAE&^�.}���3��7�BI�O��Է���l�-f�4x�|.�p9ϑkȾ�޽��H��=:����w)��U�����m]�*�����m��A�����L��W4�Z�G��\{����k��&p�
16���3&�pO�~�������HN�ʕ��m�qXȾ_3V̂�XH��́��Ʊ!��&l_�#ņ���$C�p��B)ʕ}n�U��1N$���{��o����b����@!�^��}����1kc�l5c�,{�ANr��JL���z�c�b��%j�/4�����f8Ԓ2�J������FƳj�B�H�Y��]��$L���1��s����G�>K�
���z*��鹛H���<W}�ki�4W N�u�� }��Oe���HZ:UA#�t��<􏼈��mj�ac�t�.�~�&�J��8��QAB6�t��X�vwƾ��o_{��gK�tJ��=��	%����H�I�("ҩv6@ܸ6��2��*�"�5e�K�eŭP��$$Pt�I`�@Я �,�Hnh��v2�ϩ�7v�8ӈ��I�&�^i_�-,�,���'�4 �8ԛ=+���Nܰ���}+w�B�9��MlZ�ĭ
�̞k��c�">���1Z��f��Q�3:��1�$���]�h�.�s	_v�f���A���������߈''�&ᒰLb��l,#*��!,HR�Clr��:��:�
�r*�$lBBc�$[MR����]:�~u��w"r��m��d��w�X��zd݈�P�r� ��i^|����e"�},����l�&�J;�e�c52(ew�I���(��C��^j%�����wm+h:�.)+/�O�>��������i�uD�8c�qG�2�i��V9Ijǭe�"�T�]7Й�à�H��~�2W�^�֫�+n���[͐Rx{Y�l 'i8�m��'E�Y�a2��\���r�dNM{(=��)W������hٰeg��ԒNva�@#�[tB�E"M�D��C���Dh�3��hvd�<�b�;�]���]���e�ܾ�1�ʴ�Q) �?��K��!J���Y�L!����>�^MЖ�E�1M��%cD�n~H"%��K;4ǃ��]�EE�ߣ�Bo������=tg���St;�	�O��a&�J)I�`��/�3L �t��MW��'N�!��NL�q���DC�����p<YR��R�O�3�<y�@WDA\O�b��YĹ��A�Y��G��0�EZn\%z���	��q݌}���nP&�n��$'���<.��&ؘ֗���7���"���z�O���D|��'q�c8�-���xxO�݄(-��L��/\x�y��M�\o�{�&j�����{�`�m��n��m��eЮ��}X��K;�(�En����A����#w��<eD�Y� �������;*���4ul,��;�X�A�K��0�Ҕ�.}QwG��eNw� ;�=۳-�ω�îq��.���#����e{�r�� ��噳*�
���']&�JI�һh�)�i�YF���f%����t��L4; ��Z�8Go��������'�Cq���5;�z�7n�'�ބ䅎�un�ȭi��'l,O"xڲ5�s��"����4�#��D��
���0v��\��{7��Kw���*,���e�q�0���'�k��Þ ��&�L�RG����x�u�4Taʸ��-��>��yj0����ԩ� Pgd�ۍ�!�7�m(vQe'�T������~�#X�'�7���=�
q�e�k�{����/��x��AMX:?Ź�#�Om;�����C���A�\͖b�@�ゎ�x��=�_��1��v� Gc�$��l<�i~���܅'(�"��,��:/����K���-�t�����x��=q���S&�Ym�ʼ�Z٨B�^�����%�;B*ϟ[�0L�)�I8G	�Du�٠�S�����^��d,�V�zu;�%����01��k2ϴñuO�l����گ����:F����D���Q��L䎚u�RJ{�l	KڻF�
%:&E ��<�vR{�`��J�{�\)�yd��|� )��a=I��ׯ4��+���]?^��ȎA@�)�HƩ���)��EV�r�U�ˣ�CΞI/��\"�N����&��ҁ&Q�:s�C�Ň���с�&�=��N$�l�)vQ���E��J^�'4�lA4OA�A��)7T^�[&a��	�ω�:��c���(��-�ě�B��,�E���\��u�'$�� [�������g^i�-퀗0�ɶO��6n��t�}d7�ac1�bw��q�;x3�I6��8�b����]A�qVJ[	J
�u��v�����k���PC�-��I� ���Y�ҟ�<�@B�1����R����Ypmݥ{;�35<�7���!������-4.
���3�ܭh�[(qp�����in�@j����̙����G`�. w_�p� +�Fބ�g���2���(����I�`��A���T<�]Qc�t��X:�pK�y��bP����^$B�c�v	�����F��]n_���_��n��}��y x�N"�j�R�x"��O�_�e�=Cg��f'K������c����ܑ~\�&m-E����s����-�$)G�:(�JRq�e��J���iO��)Tի �ƛGX����w�0�,�m��Lە��).P]8��p]V�:�x�'TV]HPT�[9��m�R�2V�����P�Y�!��ԥ��(
�&O%"'O�cO�9�=�*��8cP�R�LP�<e=�-�,��D����}�(,���r����tA*�^Rm�6�x�RH��޽׼��͝H
�w�n܄y�$�>�A��m�aO��a����������.>h8oA����?_�#\��I�~��]�)	��v}ksdyee������Teu�P�(��K��Ah�}46RK7ߣ��y(d��� �&���8�`���mv�Lr6����_������]n��l<��T�q���͛���d�`d�f������tX�������[Pl:��_"o��ӳ=F)eA%�;exa^����Ű��&�1�.TX�ؠ~ݓ�#�|�قUP<)E|��b5��"6��c���;�����)�}K^�f�{t:�J�I"�]��L����Q^/�݁wF¨֓�B3Ǆw�^�YB�}u��3�'������j����f��]ξ��|ؤ�uGsWR!q���V	ҳc���ĄR���m#;�����M*�-��ǚ ���$qº�
�F��]gpn��؍C;GtR�2v�*m<��s�G!x!��,?ίk�jlI%��HNv��;\��Br!�<c�t"�
8���������,�GOn���#Peq\�`$�b�,�믿qՋ�ۋWmt����F�q"�`�2Q,�KB%�xS��MeH�]��>��ʈd�m��2߀L��	��z$�g���P��`Kȇş�i���k6�>�0U4*/^z����ԅ���$���M�Oa�#�nN�U�U��řy&���o4�\����*��YD�w�%Qua����#pP�L��[�m�O�Y�����Ѳ�h�]��Y��!���A�p����KKG����{S����B`��    IDAT�$�KGd������� iGl)|] ��c�
H	|��ss�{ڋ�/��x�D�_��_������.*�d�J!�E��. M@��¨�Ã3Jhԩ�(O�4j�ʜE�I�SF(ҁ�y$6�u��MeP]W,��u�c���;�*��T�{.�w��~�]VI�2�\�'�������c���/a�щ�HB�o��Ǚ#x?���o0Y���5&�WB�	�\���U���f�%�+�/�=w�0�6?z�Zȷ)�2xt�3�z8�Ԙ�ؖYN�k�ᵋt���i�����^U���K��X��mf a���~�ڸ�u\�4``�B,���j�-D|s薌p�[��X�/�`V�(c%2�av_ �G���=V�8�5FDzN�T�w'��?�����w�kv�{f�;�����j�y�y���p>���#���Aᧃ���X.��eTD��E��9�:�DӲ�	G*R���L�Ι�͛Lޖ�X���\� �,�;y����-���D�&�gf��F�;��Ǝ ��oG����`�� ��Ӽ�Y�?9E����l��A�䓟D���%�_e��F���7�T-�Ă"�\X ��>�}
���6�#�!a��#�B�4�s|GmۮB�0"�D'��0Ϸ	G��~��ܴ��5q�QU�h���&}�4+P�6~��)�Kl���cnӊk�SJ3�>G�B��<��1�a;\�@)^��������ɕ�g�]'��<���U�Qv���>Ԝ9��L�\���\�/�
��O���ocJ��NT�2Q%Uu=�oģ��0�.���B�sP�׹���������O��^��\찂��ajj͌N�����4~�<H�d=�s�	�g��v��T�مMR�Gge�͛��ߺ�d���4�$��J���?h��G�1��8���9��e!�Z+C�*mi����|k�//m�t+��7R$�q��?������o�.8�/e�VHv��cϑ���D�,[jB���c\���%B��d���x27�k�f��@.K��жW;�y-������i~��~�;�_�F2.����c�8>OX����_Dķ@����uU��+W���pr�@�=2!&x ��M&a�DXEaqc����[R7=���
��[�IK�7��P��]��Fѻ0wU�E�>�"�P"���Lx������7����Idf�`�k��me���{���Ds��Ǜ��1���kq�<�� )a��JJ
Ֆ ��ؔ��K9�� ۰V)��>Q��i��5�6팧mZOM9�)�	G�|��#����[b�Ka��Β;$�q��s�@��_p�B� ��{g��mT��M��{~g��qU�+����"������ٵ楗^j~�7�9w�Ls�!.��e���1nM�������;�_�P=�F�RZ�xd5,�`Аi%�H(4[n%��Mfb�t�^w�Fy���<+�"G٦������~��A�
�)��Ov��ń�Clʎ�e�*�y�8j�ۨ��F��L����N��Lrw�?���/�Q�v� R-?��&\:�.+��>~�[�fQ���&�}�_�m���o�u"�A܌8�q���ֱ<�!���:�z��݃	�fe���P��]3��&'���4�;��Z%�.�l�"6L�@+���wT���A4������L/Ø��%j�EKJ�a<"�IPT`��r�+��߇R�5���_r�I��	��h�$o�����3)c���U�&���1�EU`OHoTv$VT��fcɗ`h�c]���t6�Nq?��m�+�"����l�F�P�����@4	��&�O��&��0y82��8����VHE��/�ʪ"�JY;,
ua�6`Un����\���B�����b����pM�� ��
O��]��=<�����Pږ����f9��y��h�{~k�)^:E�I��c���	�԰@��v�:7n���d�A�H���~���&=I�����8�>����]l[�p߭�ᇉ��O�$����ߙ�n~g�	�T��!����`=���{B�f�/}�K͟�髰j��j�)U��b2'g��E�O@��X��V=��F�BƮ��j��	\?�LZ	MR�,\��Rz�AK�aQ�U�M��<5	����`���e���K����U�"<)���"���Jʍ���F�A��ڈ.
��	b7��[P�;ȹ��X��<�ؓ�����n�дܼ����F�
�Zmm��� �D���529G���}�d��G����i��G�u�oG ����D�b�fg�����d���@�d��1K�9&r� ������������.�.��̹��FE�� ���țk+淶F7�A3y4|hڠjT�4LY5���7�˿��(W�����g���t����ʟ� +�� �L�<|Q5^���_݈[��;HdV��
H���-/��Eˤa)�TG��Ƒ��|�In9������l���7b:��Ѫ�IY5���z8�U�ue�mpP���EF��\~�-p�nq
6�c�g����;��c�V�3�����_�~����(Hm4H);��'�ز¹�D��k�wS�]A�ҾuZ�ƒߓ�����]��ī �`�u�ub���JKd��=�2��p����u���\�cs�R�_k(P +׆����{��V�F���� 09�G��t�xh���e؈����q����o~���_�c�qq���A�6�5��Ų��<H�0�OOAڛ�ڍ��[�����#x|�e��j<�R��Ҁ��ičmf��`a|��C7�}�^C���
�È`���;2�k]5U�:g��|5�{}{y�O-��1a܃�n�������赟z�y��w`5�X}
9�è�.ѡO4_��>�#'P�� P��p/D����6(���G�z�"ڔ6���9e9��}W�Y����9=kosks���}�2��㗸$`�8�%P��ytss�� bS�ZꣿҔ셆kcE�����n	\��~~��"���X���{U��p����}���_�|�7���)9YXx�	ʇi|ON�>�ô
O(I��w�����a��My|���nj�Έ&6#L�%-� ��XDY��I��$��۰8�;e6�RﭱU�<�sU��]V��p��?�����)�ҟ��K �n���W�h���(�#
꽷;�|��Vs�:;�鬷����0�H-�(C�L$��a$�~;���Zu�8ܯ���>����u��w���V�?k94��\�u�Wp�a� �$��Z�aw������@�IdvWNj6�2��q����E�'��}�0x���e��;� $V�l*]�����H�����?��PM� ��qg��d�ć~��~���!R��<q�,�������н�v�[��"��ܥs���{��Ï����u2����*���65.�c0+G#���]v��`������b��#�A�)ܗ��������1���*���͇/?�&���{|@�6�������_i�M<dg��*K�^E��k ��bC�������_T�H?���@��S3��`���#{��b�)��bn���'�ߎ6�B��N��}�

�Td�dr����Ϊ�bA���N�$�fq��>��ne�����]��w;�(opЄ�8��dr't+
ߏj*���_dQ�f�}_��N����� ?��U��\���w�� ��`'�x�ѧX�9�,]{�Y�}��F��&���ȱQq���1�Un����ܜ��q8.u�S�.L6Y�f�m�5T����w���Q��gP�E�wuce��>���s�.�����h�\};��MM�h�z��t�x�u.oz����E���-$��� f�	�	F4��XŶRN���BJrGP��:�ui;B�ǲ�}K�O�-�<��p�� �%r,�fUdg��%E�� ��K��Or�Eg��lЁ_ܱ���4$�b�'����ɳ�8����������'������PA5�6]P�<�-W�e�(�տ�����w����/5�=�0���i�ns
����mx��P4z�����x�y��[L��u^e,tY������1�%^+�=�W�7�X��;l:VG%�Oa�I�=v����0����܅�,6�o�.6�Hw��B�ݵ��ņ�吜\x��'>
�\�	�[o��|��y��7U�3��H3Ok�+�!�Y��	:�@��p/~���1�*��'%��g4u���Qzc��%�(�lR\�
p?��?�^"9���J&��9r��{���(�OT�V�����h�5\�؉��/G!i\������X���=��6-����d'�A�<� g�"�mo߅M��6_��d��s��<G|��;�������g�����#X�h�����Ϟ�r�zIg���de�ns�]�O��7@�7��;�P��d�9F�	*T� ��1�i�w]�$�ͥ�97C�a�f�+9w��w�xͷ�����?D�{͕7ߎ=�&��kO>�qTw/4/��F�ЅǛW�����I��+�Ҳ�~�|=<�r}�Q��)��`K9��#_~�ؾd;�T]�#L��]ڿ�uf����4�`��fgΞ�=����.g?MЦ�|�9r?�4�>{ʔ�r���w��M-.���5d60̹��@H%X���-�9!Y!�!�����l�@
�O +M�H�d&Y2�/��oTH�Ѹ^�� Sf
+wʩuwO�;��c�������=�9X���z���Dl������c�lC�<�j��z�I����:�\8�p����W�ջh"��iF��<��{������wY�tTpb�̺�=Z�/�5��l�~�4�ف�G{ԳXPt��t0WYY���=���.����WG�kWO5������o�f����,�~�
�o(���@�. ���77?�Uý $��^�a�?$D �b�D��D�tp�hwޝ_y
�ߎl\&�d>�5�c�j�g� I $�ۨ&�)b����7����{I)M��x��V����\����&:�s{4Ю<�%���m��V&�0i ~�ʂǕ����6�t�_�q3��ɰ���>�	.rV��?��4�=�W���K��|��A�����2=�Hl�Z9�\{�G4�Xs��
�p$,�<���m؞E�X[]n�.�
x���N�+�q沼ƍ��|���7���4gΝG���h+�6�Ї�����eGJan/�B � �S�6��� �������lmQP'���f��׿l���s�E.���ĳ��pI�.�sT��m�|�8	�L?ä{Q�*�St\m��nJ���J�s'WkQ?�L�������W���.�n2ď/p@z��)SS,:LN��ϡ9%O�C���M"}��]V�B�ܥ�S�a|���3\�kk2��U~=fN�Ņ�(E����}&�������泟�����[�6���	��� B�Bvj�Cl1Xm3�{�Ή�g��<DgagM{k��?�ݥ�VA�E�G=�������-������2�b�����?K�@T��ۻ�2R������M�o�m�z���^|�N�$|g1-/�Lpq��$��� ܄}��>��/M�g{����SX�fy�V�r����������j;S�̇��Cn�m��$���ڙRc�Q�;3;��qoy�mH{���P�"J��-;���
kk�})nx�?�!0�5	�3�y�{��N3Ͻ�o����ΩT�|���_��|��h��ȇ����O7���������Os��$�>�\��@Yذ�����^J���i�Y�c�P>�L�yy�F�V��MOrM�z�4����+�4��WP-8*V�����I�H��~��0��0�$��M�����	�LL��L� M���s��?�J#,}�,�g�����v��~�6�)�Q��q�¶�2�r�5��M a",AP`�9.rCb�ҫ�ؘ�;�x�^�Ն��1�Z8{f������f�+����6�D쌛��1�_�|�P�W�JI�ƺ��L��.�a�������4���������qs�҅��?�)K���9��N�U$rh�`�ץܻw
����4y��[ל�r�H��]N�e�:��Y��v�F �H�2���N�
+��v��Ύ�A�]8h����2�:�5+�N>��]�Mt��k F
>��m�ap,��F�!�2-C�6)�QM?�p!}�e��H���i	=d�ҥG��}�QD���흲s�M{�ul�_o�_191��<���� A����̘4� >��w��l��-v������2\>�'���M㷏��^�2Uܨ��h�IIfX�t���o~�y���a�d������ͧ?����s��󋁬��PTTHY�]�\ZZC6~�d%�R_ܫ��6��}�.�Ŏ�]&M��W~�n�[��`����}c�C�ud�xY4 Pz(7T�r�	�&e>1w��X��Rt�K�K��#2	����^?��>*�:~�6�)Į�E�I�f<���x�s�ɺ��31={��D���<G�92�������U�d�����I��S)T#T@�Cӈ<��A�d�ׯ��V���'3��+�wӁ+�)�&g�y
�j:�lp2�z(�Ȯ��4����Ss��cPՉ���χ}
��S��4��	w�Oq}��a
EG�>ù��(Tv����x�����U��'Sy��w86&W�pQf�� /�Q9�.&Ċ��g��U�wx�������J���~�[ï~؄e�ǧN+"�?鞶Ά�W/ܤ���izq��Wp��yn9U��ܹ�9������b*�S���A��>��>׹�q �4���B9,��M
��OX)ˎ�
��+j��7�_׿Fd�u��w;���w��v���w)�[X�B��( -+�S�ҽ���
��ߏt_��o5��՟�H���w�g>��泟�,�"�:�3���Yi���&[����f����W��|�w�������C�/����,�c� ����Z�(<=|S�*��Dd7@��(����t� �����O�j��0�:��{�lZ�@{'��.Q9�C;稫��ťK�Z��^\.�R����{���݄���Z��|���)y�0bDj��bں�॒�gE#2?����2X�L?Ӎ��`��1�o��d���H�^P.�
�
�p���&��F�ӥ�<���[���4����������'>��,��YF;�g>�S�3�<K�x�����k_��P޵���p�ɝ8�vV#��V	,�n��K��� G(l!
�,�0RN+�Y.\�D�:֡�]� �m�$���%,¡�1��I?��w��3h1D�tK;��Vit���'�^g0]�HHYB���+W��?����DH���ٳ�2qF�ћ���Qj2G)�{�":�QunX�`"�&��w+#`45b�4��J��0;;�2���"�j��>�hZ+�#Vq�8�q^TF7�za��P���7/8d��׿��X�Yo��E���v���㗛ˏ^n�g	������
[�)P��p��R�3N�P���ɲ���s����������,�c8��E���0�+	ۂ8	'�M�׶���d��=��^{f܄��i"n�Q�)�u$��]�rz�W_�
���G�>Og~d��g�,�}��mB����ۂ!�Ʌ����d�V�D�t��w��&�j���>*|ݡ�8��v�x�m�2��|A��9��*Z�=K���臨5(��G����m�[yEny��^�Ҽ���܉�mΜ?�$U\(�����Y@vl��"g8��e4q� H�+�v݀  CX��C��nvʣL�$��c���w:�a�m�LC7��N�-�
��\�ZI��E��)쫣��L��`#'9�i�d��y�[����#h"���	#8��+�ʊ[�xĖ�|u�֩��;�?,�����LC ��}6҉L�����GbšR�bX���(��qM ��8i�	��Op���8���ltU8c�EG��Nz�	l��RA8+Tٽ�^��DHzY�0�-.u�N:��}3#��*a�߃��}�[�0iZ�������U�C�t��,|8=8��I���7y����
��Xj    IDAT�:.rC��!��C��ua�<.l	��iL�l��.*��U�^p�B�
F�~�>�³�1�^�wV?���~g�Ek%�_�'"_4�X�{���@R'��}��db���pl�"��;&��q�]5"�\��u�#L���HGpC1
X����7.�
��^��Rs����:f�e����0i[�2��%��ݫW	܃��5��6�n�+��V��K�d��θ¦�R��#�mK�A��$�i�C� &L�Z�>#����p ��r���e�_Z��q'���,�O11����դ�~'Y�L�p����a2��K�N�4�b�( :ÔR�/�&�ƙf�a����zxfHH[h/QRB"ew���8X'yIw��c��v �)cn����@L���|!x����zdӱ�=H4"𐟄U��U=KZ������8��{������m0|���OyO�����:��YC�(lXa�ĻKK��X�����m�Y߇�t=hjd�̘?tG��B�;�V�P��+gE|��چդ]��n�դ��2̠����"r�qZ^/´iG�d��3��8�Ӷ���r�w�KU���bCG�n��N��@:Oܘf�uo�.;}�b�JU���z��/U3n*[��-���p%���/���Z�R���r/a�	��Z��l}[�6!�K	�o#��E��N�p�'��K�|L[�W춠VO	�+��w������\Qs�(��.K��ذ!f��V�E�F���%Y|qX��hYP��6�7�a
P�=\��%��|�a2��g:�G����gZ�1J)�u:���"��Y��$k�.�L�,���cޠ��W����S3!
J����%��ɥLN"�
ȷg�n�u��qe�UZ�;ʄ-�ηv�#��"eY�`�i��0�m�.�|��p����o�k�:�~���)�Jx���/$JIHsq���YAv�mcc:�A�G�cSnϻu��������&�����451���'�/*�A(��ul
$0(��PƢ��2'���|�V����@�q(�Mi���+v3��K#c���zR�?��F �Di�2qb,�%,�hU����gWM�K#N���$p����6�Cs��V�o�X�|�쑮a=�d{��c��)BZi����nl�(�W�X�,��9ҳ�i�U1E�,ݵ~a�¡n��>��������x���i��j�Љ�CX;e(�a���w���1=JCMAw>M��nolq��̱��tjԳ�'Bϖc�(����F �S�@2�QS��w��mc x������N�&��wڙ�a��n������_4�bf��W�C؈~OvA�;�+n}� ��2�V�!���8Y ��WsX�[���{�����"��=�h� G~a�d	�`_vİ��3L:SS��A�4�Fn�p��THr"E�%��B`G�̂E#�ȝ2���)��d\W�2��h��
f8��d���4Z��_���S��0�vD�#~I�_;]�y�߃�&�I��q3~���Ҏ|�G�3��3�0{0̃����a��a�s;,��T��)ÉK>���th���0W��\܎�����ds�kJ�1Εsa������-��o�bJ����m��gE#L�,?ϯa���-���`�t7\R��C�7��|��|�ߴ2�v�+ǍΏ�TJ���Y��˸��a���ؑ/�uzu��t"l[��~���y���3���,u��1g9�Hʹ����Zx�)�	b
I<��(g��-�A�5
!{�U:Q����<r,R�g\y0wD{!E��b�nAM�':��}Lô�����dڵ_����+o�1�=���e`/�.�}�_;ޱy�?U��I��G����w'�>��dxG�ވז%��re�>��5�V~k[�(W�Ϡ_�^�G���c�sX��O^�z�K�ޟF=Ac���؅��xo�H��sQn(2eQ���H4���,MaDz*&X8+0ht��{��q�����}0��oÛ���y��i���)��4�3�;�]��Mr3ﶺ�/!�M��@z�Nh�ǰi���m��&���@^��鵟u�poӬ�3f�i�skz���m9ĝR��#d�8�3���IC��d����`��F#	!�\��D4�J$�(o)��}Ƨ6	�t�oä��T��]��p�M��W���ƩM�g����O|ݣ��ѱ*+~�1��">M�a�4�rK��Ԅ݂*.�N��D�M/�p�c��&�yT�{/^ێ��`�m��dX���Bm���������U�:�������R;+m
���0�?j�X!nO��������V4"�c�d�t��:��+ Ȱ.����3=,^ϿM �h�_��[R�K�q2�an��i�e���|������r�wڃ駻v�e�xo�2�`ܬg�>�n\�"L5�.��i)#��/��a��3N@z�96r���Ǣ�x�E6'��<��@�XU��DP����~�DA~;*���L ��v��F�����8�[8���.W��?)��d����[��������=E��k2-��t2l	���ю���6l��μ|7M�i����H�jS���W�k�`;���	C�3����7�u���Pf��u6b��Bܨ�Ɏ$�E�6h0�D`�3zk�Α�ɱ���Z��d�0���^��*JV
ju�����6��ig������8�l��x����ey��'��8�n�緋I�ᣛ͒i��g�h�ϴ�i�y�P�o���"�j;:�v��v�=����["n�Y��2����z�q��u|���[�6�)�	��M00Cb3+���=T'�����N�<�=v�CՏ0�Gnd�/���߂�߇/�&��Ii%!Y�ao��E�(!��[�S ���n���vX��������m�:y�,q�7��Q϶>�!�V��G�L���ȡ�O�ɲ�����g���̑��0!�m=3�LCgœ���x����#���p3n�+�Kăm���%k] �*��x3�^S�u9��t��tmm>�:��C����S�m6Sx+�����(lr�0�%�U�1o�5�"��
����u��/ݵ�=�]���j��{����RQ�u����ښt�w�3���:��w�ӽ�o�����^��'�M/��O�yf�����u�7�|�N�m�i��(�rd�FNU�6�+�=tq��6Ϟ�~�#�q)w+*��A4�%���}��w':N�qA�
ʬLZ1N>�1�,�d��n/�M8��˰=C���U$�&BԈ��ie�3�(i�� O�Lw���5��l1�n#�f�C�^�(s[�3~/,�,�w�[��T�[�"�-�3=��h�w	Q(k�kg���������8��'�i����m�k��N(/~H�U�bB7"�t��7��4���q&�Aa�}�2ԋ#M�GTlaő�n(�P�ر`�Q�'Y���jx�d�0����⦿����rS#���>���du����W��nRk����n��ս~L_�|�4w�=�r�������]{X�_��^�y̝+�Pn��gR�N���v���s�9�s����#��=���e��;r���	���+G~ æ�f ��F����XAW��I��6U�tO��	�L��}ϼ|�͠{��v��3�nX��c��kZ1�gtfq��T����!������,S�����]�A�����el#�n'K��9�N;�{X�u:�_/�/;v6��t�n.E���)��Z�a�����%�%��1)2�dit���g?Op������4CI�m�*�8��^������~[���w�����n��B�=�nz�QS���aܡm|�=m� A�D�*�q#m��zؐ�K~۠��Hl�@��{�a�,�@�(S����t˴�=��'��;ߵ{���Q�v��а<���a<H�F���*�r��ylO��mV�8�]��sw	�}Az8U��fشН>1�.Az?��8;R¤\�F.�4�
r*��JU�|VT$pE�NP�u����>����'�� �1��Nʘ��]SO�q��$�k6@�x��)���5�9=�ʼ���!���E`��{���*�:nl<���ٔ��:.ZT����������Y�D��8�e}�q��x�<��?Îia舔��w�a����$d�ݢ,�u�����7M��<��١i�� N��%:��B���i<`����'h��7�=����Fan�X_��;�#ڡ?ǥ�d4���w#�����y��1�q�ݲ�-�S����l����4����9�V�o���Ŗ�%�& 3��O�5��w�hIy3��3͌���4�6N��{q9�7��=�Ю��u��ޝؓX-�o��'�_��Ʃ�qZ��H?3���薝#����V�a<W~��_Q��(ܸ���N('�����t�N��b��"��a����{�8�{�S�F�KhA����I8��Ev��V��xÌ@�q̓��o�H�6o�R?���.K棝�Y�9���43�i&�3ݴ���~��ߠ{~C�	�G��#�,�0JS�+��EpM�����0-��s�Gj��3^�=N:�kAG;0�ā<Q6���3��;9=���w�}��S��|��V "�� �[3�!a��&������=��m�fƍ~2,M����_����c�A�_�0� �]����������In��v�{ �&IE�!ːiG���"�2��Rg���F?��=~�i�g�%^v�2�::�t�]��f�דw��ά7�d���~���+k������][�`�r�
��vc�o�9�D�sߢr-2��� �"���	��0 Lҽg�n�H�8��A^��@hKy�o�밙W��w������e����g1�F��i��|ҭ�3N��N7�x�D�˷<�O~����_���y>�������6M���m�>�hX�ͭe�/��R ���o��,��[5�繁��}"�!�a��S1�vff�7]*uq��*��V��d#sT�%bg�Q�ġ�Z�N�!,)H�|�6���'#µ�v���u��}��/�&�t��L3˞��u9�{�?��|�Idlᓰ�8i��.(oG��;M/�<ZO��oq����.���"��t=�L�!0�_|q�2j���p~��'NMNL�ܾ?;7�[�A����d��
���nT����:=8�6D��T'�O;����d����ie�f�t��A;��ݰƷ��������fx�A��6����f�,����a�.�;^��K'GH�5�uI��-¶R��iK�J��S�=˯�q4q��˗C�D7ÑO��g��g�ǀ96�^���8�iT��R�%��cۛ["����H�X�@��2�X�u�1#�f>R��v�eH�gڲZ�r7��mD�!?uX���7�,������6����t>P���ii�̇�9�\ƣ0QE��巔9��FTe5�4�OR{�VD��tK_Ǎ� :Ú�&Jӳ��#��Dt�9>~j����G"���Q�C~�d����P.U�����o�MLm�r��9o��P&�������J��#'�D�
�[ �0��[��_6����&��6�,�ț�~k���A�<ـ~��1}��|�]��X����I���OiSZ�h�?P$}Y͂x�oy2/�����y������]9|�P���e\M���<(��+�&��c�l��p�X.ӊ�X�./�5n��.��E�%�w���������햍����?Ǧ�Ԉ] D�u��!d���qoทh
P�<�(��T�TZ���U�����W��_do�p H��i�/.}�g�mxJ�Ko0��ʐ����D�U�ֽ ���".˘��K�gx�f�?ː߇��yfd;�>ᇝi�ݖU�����i�S8�c���e�8D��N۴ヷ�Ep��歟����2��>6r#��S���x;�<6��M]��Np^��)��)�`Q�f�WX����A���z���DP� ��� ��A�u<�3�t��=dh��8Y��/]�M��'h�$�@�#~]��;����01F
���t}w�2LFd�d��W��-S�7�M;�%d�]6_�S�H��x�W�Ɇ�ϥ������.:���C��3���].S,HvY��rF��P>"d�K�"J�SF��AjS*��u����T�4|䏏���`���2\�#�3d�V����2e���ƫ��ib�}|�?�@ϸ�^�#�z�F<M�1�D��3T?ƕM�چ�%��h�^
�-s8�g[��_��R�0?({>~˺��k��rmm�c�����t�9>rsF T�;�F<�w�߹z�����X������De������l�D^�&a�v�m���%l�Q�K�/K��6N	[�����)��?����K���o�W+�m�,g�d"^��6qL�������o�M�Y)��d*fݨQ
��&���@H���8-�5n�G;�Ԅ0�ގ<b]�׾ѐ��5�H���لrd�H�Ȟ,.������	q�%�I������C�IA2�k)�������ٵ����+U����0����zŲ�Q��!,�����u�`�H��P5������@���42�v�>��q3�ߙv�ND����&��IEu�"N�L�ș�l��_I��-�A֩��|hĤ��*D��vVM�e�O�b��}?Y�,?��I�L�T��J�,�0x�7�z;��u�v ��@s�֭��ӳ�o��Gzf�a6sHq3N��5�\��qj�\a�+�t3�Ҋ��T!:�3s+�4TVZ�6鮛<7�0ݾ����4�=����������l�3-��hg�}���M�s4����Y�^z�G
�C�*Z�!ad�|7X]'%#��w�*��k��r����\�(��3�n	�˗/�q��Ery�3g��fKN����Ǧ�c�{���b����o����Kw�./�z������fc��Ie���R�,�4� �Ү�{�~�[Z�}�L��f�A�H�u׿��<:�a4���s����w��-"��v���j��C�j:t\mөM~�~	K���#-`�H�q2������"��uGY?��-3�}v����g7ⷡ{~m���w��w)��0��p�a]�/��/4W��aܳi�VW���D��p���ͱ����nq�����?���~��G��_���%�,�xyǁ<����*^��a�he� &�cx�]_��%���W������ ��,Wc���P�D� : rn���I';D[ j\��Y3aB�,�s�D���R��f�.A��e4>�"D�eE��R,�\&��x��	�mo�f�dC�g���ˍg�����	�b*�
�4�4GX`��A �N<H������W�� ��n'�p>y����(�G^�W
#T"s�>�O�@h������RG�R7�i�4��~�R�4^|p�扽��щ���0u!�w��X����]5����޽{���8��}�'yD+���������;��O`�i�/`5�x+���H�:G�Ѱ�N��+�Ӯ��M�	�wʑ�Y�ϲi;�v�n��Y�}�ʶ�?G6�2\)���l��)<{�>4v�o<�a�?�,_�~�a���a����=3L�~�V�~���0�G�gx�&KKKA�� ۸�4���M����#��ʠ\���3���\������A�&Y�^��ʻ����~�f�0+0�,,�!X�`�
��bC
i� $�Z���/��Eb�3�XzLO�L���-�rz��ߩzo���� �}����y�ɓ'O��Pu34x �L"TXQk�߻���5͎���#��ߒwL�$H�`�.�x�E����o���ʉ_���`9vފ��۬�DL4��X\�]&j���D�d�>��s�%����v���
8i�#��6u�q�Ӽ��p���ģb��Nެs�_p������|l�;n�e	K����i:����+�m�󷣻0�	�፧�k������T�{��M�� aS��c���}C���m�[�me�9P ���ޫA�u(�� H�)��'Ț Ͱ̿�m��qC|�9�n������ST*� �'�:�yQC*W���{`���89	��	��!�\ۜeґĖ�Ɏ�&���AÅi:�$R���    IDATz2�vQ/kk�P�(~\:��߆��EF�"��n�7�#n�O�7<g��oې��?�1L=wҏ��<�Qka�ߦ���7q�l/��>�&7+��ܡ���S�o�C�
�>*t+p*�%\��@Pb�w��!��iZ 9@ƿW�Z����P���x	e{�Y_�,�'��[F3���~�%�Pm�{��y9W�v.9�:)p�D9U����(�6!l�Q9�Sۦ�G�-�Z�KyN���j�j�B$EK��N�����Z]�1�i `���m�E>�Ƚu�%Hb�q�V�k���i�!�5�_8�����e�[{��o���0�ۦ�U�
�3�7J�M��76̌:n�����FG�6�  �#�f���qr�'; ɢlP4>=x�˯?�͸��K?�I���f���2,�R�5�tƱlo+ST�N6k��v�q�[˴_W�hsnwNE6]�Q��Xyӄ�Q��<�P��5�Z.0�3.��SG�����00�I�n�lk�}/�j�*�eX3��2M�3N3�f�2���WK;Ju�R�m�E�����qk,�s[s��V;�~�(Cx����Jg#�a�9u�����lp��Ώ�>R������Ęqrk	�щ����!u<�y�1�O��wn��Pc*��w�+����Ǫ�@�Ͻ��e�Cekr@��`��D��Y���e�9�%��!acT&�d�z3g�trx5V��~�3^�H���g�n<ȸ|�T���n>�4�t�6�ȷ7FJ~���c��Lo�$l;�D�O�6���v�p�%w���/����n�_�At�K W�����M�I��?ٰ��6<1��4��;�3�j�(_��n��������-����׶3��29Zpb��1�5�#՟���N�=Y�?i1.��].G*+����!���O<W_E�����r�b-�J@I�v���8I�����('�ǯ����r��\l'��Єg���g�a�m��M8�d�(�8�.����~�4��Ҁ���靃({[�b�߈pX�m�o����Y�ܖ�����?�t�؉ٹ�Yv1T1E�XyS��_]V�J�x	�l�a�峍���3N�D�@�pަI@gj�!�s6��oE���t�k���b>!�P��E�qɸ�7*�������~���/y�;ʙS'�[�r��yzv�����Y��@T�O����g~�_��7��a���M�P�,��n�G���h��o��!���O��0�j��/jh�;@���y�j�5o��EZe)]ԧ��߰�'���y���QRF�O�L���V��h]��-#ܶ�0?yة��[��[F��z�_&Q�}hKX��s�f�gʥK��&g&O��j �ȡ1>: �uM��8�g<��7�n�����_$|!NB�� T�@�1qR�0��.D8p�]������#,�,/�I6ʻ�����|gy�����F�=���A\�f�7р�H���n��ɢ�n��Un����������/�ŏ��ÃC���7ʇ>h�)�W�];Kg����m��Ω(C쀭�&<~���o�����4��m�$Ќ��ɷ����;4�q�i-#�}�Kt��Uƈ��Y��ǟ}7[aڬRm-R� 㤳����O�M���È�@�{��g����������S�P�Վ!�3>P�a�	����9���4���c�@ME���㮬,w&4-n�],�������a�������3g�F��;������t���Ъ%AL�Z/�+Kс�ۨ�P��n�@�̗>U�㻾���o����� � ���#߸G�vKW����au��m!Ǉ�����f��ſ�ᨶ������e�q�m$����5��6]0�x�N\>F�L:��q�dX�M�d��D,A�F���x�@_�@{re�3�xß}7�!��t�{p�Ņ��Y�=������К�͜��I'	 l��?�N���̣Ǹ��N��n4�yBt0�^�hSG�8-v�&�,©����ʷ������?/���x��ܭr��edt���=�텐�Gǆ�2HPk�ۏN{��^��^,m�#��gv~�0�5������|�,΁L��H9�O�˶�	�KOo�t���:�Ǫq���F�He%����� ���[M�"�R�O��~�8M��	� P��6��f�13��X��ۺ��������3o�c>�x�˚Ag㼑`�웸U2o��ͱ����S���.]�|�����@T�Q����h�g:��8��ЩJ@����j琯�6���R.5L��w�ÕZ�u�G?2v�d�!qjz�<:V~�����)O<�tp��7����H�mM�P�����Kޜ���\j)�ss�29�k
��7�5���|��`5�P)s� X���A��o� � ެC���.�;�sQ�
\��=���6���X�
�J�D�m����a�*�/�z���:�6c���-F��9�tF^)R���0��d;���\Gn�D�ށ�m�d�Y��o�6'
��,�щ���-��s�6�����Z'^YjT������26"]�gC�?߻�6�3����8	@�ã#\?����g�BY�+r�U�?�ߖ�]�QN�8VZ�}{�vi��0�0�K�V�a�ٰ�_(�䱶��|�P������ksL {�3��.R��/����\Y�X(0� |����2�\F��n�3���G)s+(f�DR.�dm�KN�K��n£����L�y���4��n�_~�G>7t��诬��E�)�����D�:<dO�o�V�`�����'�li�966�+[V ��a$��?6��0g����{�7��"O=q�n~��Ov�9�=9�0����|��{��<������-�mO<^nܺNf=eim��,VʁC�M$ N�,K�a�Ņ��K�(tn�[Y[(K���Y����UeN:bIԍ��2�����C�-��(�T�C�O=���V,��j�=5����U�Xu�f�颭�X%��7�%����;Z������:���¹�o]���|�=�UV�6���89�J�T���F����W��{n~�d�}:�p�9�z��Iy��-f�}KK�C�����:�A�Z�d6���iX9�9��Xc�L�O���ٔ��{�,O��K��dp�<8Q��뾮��/�<��G���g�0�v��,hJL;=WO�w��6���ѰeĔ����؊&+�p}k�q�hKBd�x^ڵ��qtx�\�~���^,��?�n�zQA�]�ss�,a
{���r���N�=S�H�� "Oߌm�vO�)`[�.`%<������?k"$�vǈ|:�)v4�J�%��iį.�,�wı}�/�ŏ�0vt��2=3]&����9��훸�v���n�i��GZ;42�422�b���BD %"�UW�X��y�٨�/|�;�6y�="�'�bz�6��.��:9�����ȷ�3�;�-���o��������������-?�3��,b�8��X� ��eF��!؇ö�K�=�\�|�}�K+�c7������Pk�](]}��@��� K�uu��i�Q�G0{EDi�_�n[e�`wz��8p�<��g�����K��G?�2wg	9��ϔ2��0~`��۩6�Y��.m��+�.,Y�#����n��� M�&bL����o�ո��$�:�1L���HO��h|7�PW9���O�f4#��#A�L�[�-�����RYX\ w�V���ӲN.O���M����H�nB4��f�jn߹Ӻ35}�ƍ��rC+r/�� ���fx�U ��o��Wxm�������p�$�*/ S_*�O"�_���]�*_�~��'�SSwB[6�X�4 �A\���OȡoܜD.$��M:�~�et��������#�aq�E�ۓUMj��6S�5F��h��p9��q./��[�7^���O�x����R����-�{���0�.�=r��KmW���.᫖�F��$NF��2��h3����w�%<+�Ubn��;␮7sI��̞B��S|����5?q�S���1D�eĿ���-\e`��훸=f���2����JЃ�]#�肆�v��o�Gm�@�����{��ߘV����,�I�����|L��&��u��ˋ��������Q~���Us3�����7�!�jiK$r
��B�=��$���opS�2��YB�1��-#��b��Vy�«�7��[7��;�b�I����cTa�����9D�6��V1f�A�(;�F��0������ղ�:�:�U��-�*O<�X�uy�������k�X�Dg6V��c����d����
c���C��ֶ�D�7�Bh�1���vʻD�N���1$�T,��U;��Tg��ša�j673#�p\X�Z��T��"���M�� �1�a��X�`p�P>0q`��x"=�F�ƭ��׎s�`<�Kx�W6�����ɶl��^�t���2���P)���G�G�?�����_�;0Y�2�0
�WK����y�g��z�.�0s��M��S�����r����g�`���j��A�GN+g>����zp�"2�P\��*Q�W��[�f�p���z���/�wXb"�B]��Ï���vy�3/R�Fy�˞(�=|��?���eq���m�
m�� #��=ȩNb-��C��X!:쿙K���?q��t�߻�3V3O񞋌���nA�Ue�$甌Eݧ����R|:�;{߉�eD��ܛ�n�T��׹.Qi+nQ�S�d��eG��"�w�P�m`d��x�c��)�����5�~�cE�w/�2� �����d��gx������?�? f�@��Qg�͋9�u4#/��b9u��;dr�&����1uy�u�Y+g�?!v����˅K��(�O.�xf3Z��c�)�G�����2�`z��5��AȜ�;`��i'<|�H9x� ��iĊR.�|s�Vy���Pa.�˯�/�#c����������}���⫗�X�̈́a���KBU&L��qx�/ A�w=����t�:V#�s�?�m>Y�6����iS���$�N��By��-DV�;W������ު�웸X�:�����/�e����X�7�l�oh��B�S�t�5N ���ݶ�̼���G�SV�!�"�f��o��o.?�/�r���a]q������/?V�#O<B��GE�9oay5�mD��r�ܩ�>��Ǣ�}h�z��2<1T�f�ʵ;�����L�0�Va� ��"dx8uϘ�౔�v3�숽ě`Yd����-�
��a���4��b���+/����+o��'ʍk7�s/|�|�S_�X�E���/�Ͻ�j�7��
QJbvBg/'ﺀ+p��Y���[�k��F'yg~7��<��bĕF����S�ڕ�exd ����o�N��܍�����}7�ބ��J9�;̳S���.��u'��w���-� 8��O�]�3��qI.���څ�P*`�_#8�.�a��y��5�������-?�S�c9}�L�]���/UKw�߄p�˷~�{���$\e	�y�ܞ�Ew�����O
���W�^-c��T-��*C��f�E!���xU�ܕ	%�a��D�b�Z�Ů������ˍ��W4��3���s��XC�^@C32�.~1g�0��r������k����˷�?*���(]��_��/ï�p��MD�U�(�rw7��*�T;\Z�U"6<ݽ1��ɰL~d��M��ծ��l嶱
�@Z#�7��p^�=�&j����o���m�u�:+g,��ғ&�*ہD\i�
�X�%�jl���w�w Jw2i��8��W>�������1;����So��������Ν�ஊ+��.O��_+�,��6cf��<R�_z�|�._��_ZN�=�n�r��Zƒ����X?�ݴ`gҶ$:�256*m���+�s[S����W/�R�#b<x�zpN�A�d	�����X�^�a�}��Ce��hy��G��+����}ٺ]y������WED]߂q�F���>������X��I�:j�n9z^	cGфa��w �?�I|���m��;�o<�����̟��(�7�k��˪��ʚUP���/��6��Z��)�"	����l��y��WƬ�ĩX���� ��-�͆[�Z������[c^�E~��t�ޙ�]�?�H�ٟ�9v�� b`>	\e�ThZ��uџB�mT|�Ja�ň�z�tY�/>�e
N��?��+�g�8P��h([� �8�4;U�f�Y�\@��}>;��b�s۶�v4�:t�@���̡j��Q�Ⅸ3\����1�tN��[��}��K��.^//��jy��g�[������gXI=T>��O2�`'s{��y{��-����t�G�#�쌎����a�)q��I?���[���u�|�g���M�>DA��<MWEv+������������=�~��{A�p���k�*6+�j��k���+�	���֤k� ��d�K���۷��%L B_.g��aLy�o9��YA��s?����w��!m>�˹�t�o#W�e=�E.���_(G���G�-��w��/}�Xyۃ��o��8�(I�a���e}���$
6F�~�w�GЉ�$ƦD�nԌ�c�Ľg��5�Zc.��?:!b�,FC���e|x<��r���#��&-/~����|�|�}e9���2s{�P�o��o*�G���~��R���PAv��w��a]q �	7��O���N�8#��:�}$d]�[G����b�:0`+Yı�۷�o΀���.B��7D�KU��d	�sL����B^db��r/�  ��p3��s�L�| f.����I`{ԣ����1쒧r�:6���� �����/��������{�ɐ[����L;��=qd���xp���-�k�A�}��b5t����d�B��;��q#G�չ����$�z
���t��Q�z�\���jR�Ս���[pDH$d��6an_��m���i������c|��Վ,-!����Ĵuji�ej�/�_R.�r���G?X�|����S��O~�S�U��Uϔ?��?�6C-�փz�Is���Ĩ�p��ĭ_f�?Zx�G[�h2N�#�#.�Y@��������[�$۲�TN"�A�>6::�r�F��Hq�?�&n6�`������O�b����L(?��c�r�>I�����!>�����@�u���L�o�3�^���Պ���0;�����?F�mv{��L,���E�$�~G��ߚ���x觗]���?�ɏ K��'Y49|�@�'��׮�ZΣ��B����h:�Zȥ=|G⎉2V���D�	�
��Tn�Q�:���T�F�t�W�C3`۴� �5��W!�j\�8x�H�9}��_%���G�'���v�|�g��o�j��+���[~�W~����kl��d`n��U�J�6��u�Z�^��vV����7���o��_~'�7��;�x��0�W�b��b�żzt��	�n��=҉�S[ �" +�۳�aL�P=���q	 �l���#˩u�'����_�k~�|���N����k�c�OS���,����Q����I�\�}��[AE�_dw���#e�=SfYJ�ӟ.g:G--f��3�0�2�tKM��0�V�vG�L�Xu�@�j�f�PB���E�=t2H��U]7D��5aD�m;�E]{����z���՛�ባ�ߔu}��By�'�j��+�˥[��S_�ty��"�L�Ǟz�L�b|����u]�đP�x:�Z�V���Q>J���:F<�4q�'d�w5N�%��ȗ��v$�q���/��'9�D���k�9������[\��o�^n�7U�"�޺y+��yn/^���>1b�3r�g������o��t���w'��oôs���lC��
_pRc���7?���=��&v�L`x�b������7��FO3+!_�6#����it���aӱ�A�,�}s�:K����Ct$�g�<
D�K���d$aS��"R�7ce>�!\�Y���4��h��1;��h�cP�ҋ͈�wX=�0���{ј�o���g�8Sg��	?�Fe�<�����#�ș���W^/��,�=��5�[�X�D���?��r��l��	�čL��u�W	N&�V\    IDAT�5�6�Q�.��m�fX����;eV%@�;g���˗#^�/ 3Eq��p�pwS�w������\�p��%+t�����/z{칷�I�6R���x�w?�0�����_~����0���-@��D��?�c��qrj2��89GP�V�я�fQ�E!h���?�C�Ҟr��1�Z(w�$��r��A�#,��D|9x�P醐{GF�h^*�;FG&�ɓg!^�*�:#�;���\�[�a�{��G/�^������},"m"֬l����$WRG �^��[,r��&Y�Y�.e��>��'��s.�u��W_cԂ����uy拟.GQ}R�O�Px�q�.��q�c�B?���;:�,��W��N���V9z�(�EN^��/qc�?�C'�7����7F���g?�kiq4ڞN���\���#nd��A�lN�+�;���4i�|"��������-Ӹ+��~��2t���V`q��I���Q��}��˷Xf�x����g�!��X��d�\�q�̈�bM���G@\l&�hx)�S���hvy�6jŀ���E	C��K�۶�"$�.Dq��X�uH�� ��01�\ԛ$��!������X�y�v�ڭ�V�5aPn1�@?~��!�$��#���Yn_��_U._�T.�!���&���o��7�g<ã=��t�#]�J|�<	%NƋ| F���T�:E�d����B,��ٴ��+3��YT���g����Z�*���u�!�Ǭv����r��;7[�[	eE	@B�Qx���r����$�rFc����� �+������ �mZj:�?��B��;W�����2���Y��W�m�%�vn"�ݙ�]&O`�U�7��?W��6�c_�X��Q���e��]6lI�c�^�w!E�E?n�\i��6:f�����Uİ�C�?N�<"^L")�{�:��l���8�~���:�?�mN��S���#�SNkh�^���EwD��0�]���<�m����O�-�?�jy��Ǣ/������>\.��>�N���d5���p�zhgM1�&����#���c�S�m��4pD���G�w>�|�I��㝂6�p�g�OcW�[}23���c/��!n�cо��/qo��3����N�!P*��v�>���h����x=4��S��߫nٻk�#�W��۞/ �ܷ��&�9����uo�6պ�)�����(7��pX΍����h�����by��M6,�DgfC��u�x8)5�6D�2�\f�c/m�u�����R��3�l	T� �b�Z�,��a�����26Z;>\
z��ʜ���H�7�!g֕M:���vC5g�l��WY���|ײ�0���s�4���S�~�Xz��'Y�����0;�PR��a4H�1� (���	{�xI�gr^�����q���㛯����3/�\��"©�y���,���X�][�A)jX�#G��[�o�k �����t���[�l��l`>��o�R���@nz����\y��u:���'d}��锹gf���6�Ͻ�\y�[L�yЉO�Yw�?y�:z�u����6�]H!Zx���7���Sw�%�E�ι<h%P�u#���mq��ۦ�׽�N�5�b�[[�艇, S��c)XB���g�0sa�sw���*���F���~�3&���7nÙQM>����/>W�����(���-o������ ���%�L���n�$>�đ��N���t7��wtWI��Y��������%p�7��f���/���]0D�n !8e!r\��>�����Y���A��葮H���a>�݁c��{w���4WN$�y��?��1�΂��� �E������ٍ��r��q|�\�v�vk5�-ƙΔnV��[;<kw-׆W��axU�F$�Sk�d��VUY��w��]C�-��~�#~��
c�oa3�}�ڑW�A�����!Z�9^ �l���̅!��FY]� 
},���"������?t��ȞNl�~�����ʱ#tX����a�_x�,#�n9v��:7J�'��x��,wkP2�n<ݝί꤁��q;]0�z3�LI7�0��`�V3i5�[r�}7̢zƞeo��67��>����Y�$���H��Vmf%���[@e�0��7"��c�ݡ��}�� l{���c�c�6G�D�Z�M�sp����E������W��Ȳ9m���n�m�8�V����О���
OèM�z�,t��J����Cs��݇ȱj$MV��w�j�$�i<�P�B;W���.�ۑ���@n���!p�U/��]QN��v!�r|c��W;����=p���U^�z�<p�2�>�.gΝ)/>�
p���.q�L�^��w��q�2xԏt�eG�%n�u(P��x��X
�v�&̛���8��� ��V����`�CSiD�&r��lx����-�i�f�ɰ�6���ÕFw��)�W�D]l����! 츽K��6.��v'�g�2l_G�
\}���D�]I7�,�s!(6 �Hp����.Z}��Y^nn�`�ǈ�[M���S��'�Jؚ�
�8�U��Yͅ�d��=�
�|�����ܱ1��~h;89�Ot���тY!*�W(YWG�뷯���0�������?�YT�'����?�hy���uz�2���`OHGb�9;p��(D�S���H�������0]�c�3m��N<��ϑ݉��u�rY|ۦ�f�o�:`x�Xo��"�8�G.)wH�0�h��٘l���>�	Wߦ_5ߑJ�G��f_���|��} T 	�:�\Ἶe8�;cf�/_�T>�z=��<�!��!��%���&���e&|څT��#R�c0"'��p�t�y�ܶ�Q��<�xp�?^F��YJg`�G�uT��>�B�tT5-��:�|�!��i�o~#�@ �w�ࢢ��v\.��C���6w��E�+}���qt����:o�j�l�]��h{��� #�b�6d&��th�r��"d��|�&���?���0��3�;o�+�G:��,l�.�<�;a�{�Ľ5>�օ9�G�HU�>{�lp	�J�VT��I���ݰ�w�4��yd���%}�;�*N\u3�gjP�����nZ�V7%�m��+7/ý��Q-(�o1�rgMplf��A���JH���q�25�A�ѷ�q^q!�4���=,ǐy��4��6Z�iF�ؒ_���"C��^B4�*�ؽ�́?����+������?�8���7&�pl��HΈC��I�ѻ1�y�P/։�L��f&cdz�	�G­xPmWc����8�@Bd
w;�m��4�M�\G��1މ?�~���<���w�'��`N7n�(ׯ_�<�0m����֤M�Nw3��~��Ĳ�:���6�G��_�5_"����a�����l@�ec}g\�(��g޾M�oӛ��l�yNc�t�/���"�+;4�EC��>ȉ��h\	�=ѻ"�%�"�ݦ��/bҪ�����D
�3�4xB}�\m27:R���A�X>zQ�ͳ���(ps�N������,�ϗe&zn4�]��7�Nx�\���\#��ɽa�n�v��x��v�∓N���qք+pp��8�l(�n��,@qM�.'��{��r,�,���@9�~MՈ�OpjzM2(�(�+L+!JĆ��čp3N�ķaMB׿�.���r|�0+N�\��o�kq�'��Mܾ�{dd����JX�C� pO���$D`���� �1�$N���o�y���Y9L�f�D�q�?:ĮA�'E�(nܐ���{Y�^�xV�!�qs�c)g�CE�ї�3�`O����zƙ��c��Ǆ2���ȔWm���pkb|{k�D��Ԋ�n\��o�;�e���[lfq�>��V*>m�
���/W��W���s�F���U���n�	�~��aeՑ�c.^�j?��N�+����g���2�<�����A
�g�w�@q3�/����@ša�G��4]������m{9q,�:u�T���{i�c��j���9����z�������+fu�*���0%��}��Qy�6�FAST�Y}�f+�8�q�O��?�w �]�r�U4��4��TF�)�&�r� L�9�A���������tp��FP+�R���P��^ۼ�������7V�'����y��B�j)���W��[#�qW���.a�@Ⱥn��J����AڸH��Ȋ�ת0t��o'���K��l��r/b�O����w�	��)�8���q���\�!�	&�m���<&�k�Kݿ#��*�����r��U��N<�����������y�o'�jJ\\�a�8����\�|o��K��?��	A���}c}��	E�V\�'����9[Q������&�鯘��cK����	�R���y��7~�7F\'fZ�b[��Y74x����Јx �;h���%u-����ۊ�W�U���2��gr�(rl�x |yq�+hK}�n���y�bF���ys.�*"��q���M�Uֹ;`$����?�g�8uJ�S�{#sR^���4|��4u�j�7��G���+�ۮ��Ƹ��fp�I��y�|���娊���8��5 a�?2���1G��y���y+׌�� P[���3N�Ź����:�S:��p6:�/��s{�#��A[��pP�w�F�ج�o��ț=׼m���trg��v��3�~�y�~?��?�&�r��T��c\ۆ�8D��]PT�c%���fPNh'��Ғ�1�+Vݳ8��"����������*>*�ɟ�I$P�Ze"��i�'��lr�D�N�ـ�	)k=�YU�M�u��Q�l�v�Q��<�r����HG�u���$J�u܍�h��q�͵'Y��V�v�q�Ѓln���	�g��=|XUj�E�N�n0��¾�$��'��ﬣ�L��淿���xQ�I��n��s���n��#�� en�ەH� �;w.& %V(�+���ƷWJ|>��Cg��w>~擝i����8Z�2�zw�(Y��Z�T�\5'KL��#�0��H�dzp��,�q&6��P!����I�N��&MZ���Z�8�n�Jc����R��M�/v��:r�\���p^�#��i��m_�Q�\]QMXȤ�A�U|����Ś��C9w2ML7�f�G�!����q��.�{�n�x����ʴ�ru�M\�N(�����,]�:����?��<�-�ģ8�F�W'N�W�YY9�'q�W,	��{�u~�=NK��iNG:�p��Hl���P��F�[i+o>w�7��Q:�����mfNN�F�4z�ɤN@̡�0m�Jױـ�(�NH�[���RX�!bH\N���ejy�^L���L�B�*���N��@�=e!;�!K����|X���à�3��Lԝ3�T����-�I$�@��� `^�e������ꤒX�W��"�"�(/�����­w���z����3�Y)�=[����Z7�x�z�>|s�Q�Y��Gv�0��xO:˭e���������^��ү���_����_|8��c�$Y������so(s�����X	���y��`1�&qZ)�~f�[ �[?�C��o��(��<-[?˲�ۡ���1���l�8"ӎb����V.7�"�i�N�\Sa�d��O�S�b���y�rtȝrn�M��z�5S���ud@�ww�
O�S����@�:����/��w����\����E����aX�9��QW���>N��n�]�2X�{�$H�`'1^��cY�7n�e=�m]~�n�l��q�[�ąODʼ���z��g+�k&n��/qCT��=��+ �E58�N-q���:Z��z��)4�I�@[a'8"N�	|+l��=T=��~"���G�F�-|���f��,�Y���*�}7Co7'��[f�N�����nsvv�{�	ey�O�b	_]�`����u����6���#����G�*��?Z�Cp4�L�>��P[ro��͞�����"g�wqb�&�1�g�B���M����e�	���o%2`����A�5���vb�(&���ݎ*t:�2���ު��B�k'S����g�b s���w�GM�@}5,S���/�c�+�k�aֺ*G�]�`�1�-�"N`!>��Aa�u���l�����8�m<�|�ʫy��+3�m1��p7Y�P��5_�n�a����;	�k�8o��K�QqKN�!�H �>}:z��)FH���f/mt�SbO��~�%�$~�q��ϕ�U�\�>`y�V��.����\N�,�R+����'��7���se�x./ /[?�thR�Gʦ�%�;_�v�{�E�И�?���x�?]��A��뗣���Qb�D��f��z�͵�Ç9��)R�i<�1��-WƔ��e�����eX�ɷaͧɸ�o�.���ā�^���辐KV�K�Q�GU]�d=��H@Y�l�a�����<����	��ph���&׶�Vݰ�D��䁚�# D���3��.o+�:s21g8^�Su�+��������G_<ZEқ�h�y��n��.��Ṳk�!` 'KgX����3~�;��rP&��(y���]�(�y��+�^deG��N_�92���d��K<>�ϝO�~xêz����m&m�E�p~q-���0d����y+������}���E&�[]�2�D�+��R�\����S.gX:�� ʷ��	x�D�.���;���VW��"�H�ޭ~���,u�M����g9n8Xw�(a�Ѣ� @��{<�b�5��b�&�t�\�6L"�5�zA�Q�=�ؖlF?>���m+~A�ؙ&�u��l~7��mÞ�	3��y��n�D�@hgU1��&�Z��<��O�۰��o��x��w��v�^g�O�Ȉ�J��7o��u�4����CA�
��occ�k����܃�m�Z�X"a:���V<���o�.�ˆF��aX	T�'�;[WÀ��f��#�s�w/gs��42G5$�&r3`�p�|2�A�ڊ���"W,��rc�F�v�R���S����R� 	�oN;.�HL�сb'�F������>FM�*ڪ8$��D�-;Dc�S�c����D�;��>�%l�.�!vۤ��Q,�yZT��L���8��w*,�m?�Lox���������E5�?�$�[gq���S����^�
�{�|~X��KX)�Z�"B6��It6�	lM���8	�f��'�1<�c:;�gS�>�9�:�f��$�-��b7��� nI���)��H#�-�eN�0$A�Fs�N�S�\��9�\�O⋣�E '���{o�[�!Ĝ�R�����v]��w�0k��l�)���W���D��^�M���Y�FW	��2�ϲ�S��Y�5�߸鯟�ű�r�����/�\��IA����&xwo(�I�wP����o�c���D�E+?�L];�l��|��~� ��H��wܐE<�~�o��GU|:;�y&p��m�vܞ]�VŹ�����B�ƸA���w��B�#�ߛgٚ3˥+���{vӭ��h趰�Hul�u�o�=���(�<L�B����M'R�o2śq�pk���ٮ�.��M�c Nʹ�U�~w)����M��w:��N���?��۸Q�J�y��0���6���#������K��~K�)��s)\��^Ugeu�;��^����|���  �K`�n"�o��!V��5���tTB���f�26;;���7�-��$j��˵���Ԍ���._|���q+Xj_�6����кHt��؎h/�t�M ���	kM��#��6]�G���t�j&.5ϝ��"y).9Q�d+��S2��Q&d�M|BcB�_�3jM�IPg�a}��䍸Q�[�i���v` ��;
�ߑy*UF�u#ORo�Zܥ�W�>v��'Y1��yf4s��������/�8޹�H}�9��<�z��>����:�[��I����� ������Z1���ɫe��+�`♧H�\ì������[�٥�ȗ�9ْ�E���V]=��fh`\���V��i�>Q9�@��m���T���$���    IDAT�"����ݕ/�ԲjyvFj�����3�n���t�[�D����%6?ce��Cq��*A�&βl�0�O�ee}2ܸ:�3ν�#R��L�x:w�\�H[�np�ihMjo�{��7q�����0�b���$UoVІ����a�K�>��۴�o����P߆�N�o��S� B@��<{��=��{��oZ{���q%�2�r��3�l'����u�'W��X'�Y7�u��t��p�-�'��L�w��v�$�����2?���B�pÎ�p�5	.�aF�2��pgQG1��^�|�/�U�f�(3PP��QF�%�������W�%2�2'���O��������7q�8�ծUO"M�{��)sأG��s[)+�pW�[D�X	�C �gw��&Adߵ�TM�6-ADi��v/�-�܍���v��S��)$��DU�79��H�WC��Nc�j�U$��q�G���(/�MK��H�[��55���!
UTO�Dr���h��1�w��ζC�~7;����8v{r�ۣ�U� �э���1ɚQ�_�"t�*a6�%Y�,�r����V}��$ئ_��|�Gɜ��ܪ��ѷ�M�u4���o�^\��(�C�	���/�D-a+s'w � �o�M��?	�8����Ir����␳j��n�r��+���k�D�ܵ���G��C:9v��1ALJ�Sw���QY�C����ݠ��YO�p0~�)��=�&�7;�u�~�����L+����s3�� ��vb�D��&N;��\��E4���
�if�Ik���wʾ�\kgX�1��w>����mJ����V�Z�Y)v:*G~&?��{��ƀ�~������_�P�������d�<��y��	�b�E�Kb�m�D��x��ƿ���U>�W��p��� !"_���6/Ü���e�,W���Q}�#�>��f��s���zsø��DE���E)�H���@fT����xUd�|L˓�Z��W-G¢^�����|��+ض�d|�ʡ�ġs��\���� A{є����p���&%�!�#����E�Ο,7:����i���1�D�w:q��̷�X��K'M�kGcӰf�>�~��C6���kH�v�H`��ʲw9|˥tV2��W����4�_��6,���@棿�+7��~����y���>=����U�7/���?��D�dS���qm��[��p	X�K:��+�'�y8��m��g;��v���!�ng;v��1���,+�Q�R�ɽ%p�77�E���r��Wr��?���f����[<6?tڴ��Y^�C������u��~7��ͷ\[KԊ��,�!��h%�f���=���S��(�W�M��%2�<��F�Vfˊ4ߙ�~"/��_��~"!�d�v���Mf�٣}�]5�ҙ^"�N$��[���o��+�FԈ�h��m�ۘp�屢���+��}&�RUM�,����������`h�rl-?�_������s�K��~��X/��-A�]�-�[��ϕW���Nr���Op ��\[!W7�OmCe���#-��?�����j���n�f���uζK�rleo��S�sc�Z5{�]�Y���*��j�d�Y��w�V8e��n�nW1��(���)����Ĭ��-W��4^e�#�V�{�ز�鎥�NW�u�[�,����=q6�)zYO�ȩ^	pv�3OãL���.�f�Y��w�hr�L��������,/�3o9��6���ܹs���[1J-1�t2��1^���M���N�e5����n�5ͽ�-O�[)�]m>�0�Z�Ú���;T���g7�b���.���_*/��*�a�,CC�/w4^;\�T��𽡂�6$A[7+-&�"�2�� �����K����v���3n�nۃg>��gم�7�8����K��#`Clkh����.�Or��&�؟�;�!$8��;�1����r~��s�l�8u9������K88��
�-�ԌE$�F���s�\<`��U\,aBL�`My���E���b8�\��hÃF�7u��c���\�D'N��� �}�U��]�p�a�v�-���(ko9F�=��R9�om����x�!���X�c�1x6v�{r����N{7)o 3��^�������1�|�g�~�ֺ��{	�I�,'�^s;g�p�U�7׻p�}[	Z&�5О��T���r��8x�����aE�N��X�r�2�k������I����	�㷆:�����L˰<{�K/��<1�ɵU	Z4�����M����	RYo��\[�S��H��>�qƣܻ\v�fź�f�ߺ���ٮm����B��m]2��|"���6��e[|r4���G�˷��0�-G����ə։�pS���6��䕗^�ޗaL�N�~ۮp��|u��0}�c[��ߝ��_�8z淿~���Xݶ���r�6�=�3ܓ~����B���D���_��awۼS�(&d'�2�B��ߍh�m\�v��#�Ry�2_����/��/���8	`��=�Wm��3��2p{;�� �E��;ʈ땜��z��w
�a�躇�X���?7{�k�	gi=K}lK����lN��u֥�}g�JX�q���|��R��[<���N$,�>5�e:1t/h=�MR���Q�y[⒬��/E��<�����N�td�"�c�C�GM��v�K��߸�O2ڍk������%n�P��`*�-�{O훸ٟ�α
}K�vEP��u�vk6Ԋ&��2�͸�N.p�F'�/�Ti��s�e���O~�\�u3��L<�X�������d�"����I�|:!���p�SRo,�t���{���#�7=j���){Kt�:�V��N���#��X��K�Pm�Y�z���]�6��0|n��_Hnz��x5����M=����]:�_l��N�W^y�56>#��+w�"��;eG��~3��t@�eܨC4h'e3<}Mo3,���0m�Th�=����2��.8�n�Ľ���Ĩ}59�e8t�w�}q��L���������x	�Ls�w�y�9��〕C̡��|����=� [�Z�fc������AҰ�`�T�D���x+'ֻ3Q/����0��T���\#�?�+���X4o �>����|���}���5�a�>�\�ݖ�a�����������h��Mp�J���q<���B>|�6�w��8�[�<C��#��y��� G��Wn�Gy�|���C*�@���H�ȗ.��B��'YՇ�&������%!�q�/��;��R�b�����A�*-EوB4���7q�goO���S9۞%�;	���o%0 Aq�)����Fuz��q�&���;�gy�^�I˕s��O�4G���H���V�>��߁����|Cq�R"ϕ� (&O��}{z��E08b�]�)�.��o�^�8*�KW���[ԩH��8	�k�$s��^,$�����x98t�Ӟ����f�� �ND��#��ƅ$T�mgKD7q�p�~ �+�߆!��;�+^�Eы%8��3Uf9�����}��0�]�c�7�R;�"���F#����������C�Y7�w�=������f;$b���y�����g���O�	T���n��7O�Y!�}�.C��+	׳��������9i>V>VOi���l`�8���z����v?�@X�Vgի삯r.܊�u�
��96ػK[�8e���&ǌ�,�jb��K�%4��j�Zը��B�X��ߘ���dM��o<S�s�u!8*�-�?	���QB���7\��	d�M�!(�@I�5pD`!l��`v��-�A�V��?d����/`�_F��h�J�:�=��o��Y[\/�7�b��ǅT�}�����O�K��+Ƞ�Ipz��Й�E�#��7�	{��k��u�����;��|d���z�37pB̂a�۶�J��-�l!w�W4�$w�}s��ծNq�V���F9��7��YBO.�\�4�o��N�V��is��pe�D��/��b������K�CTpqb�[\��� �fń�yVV9�b��� ;��zk�y�X����ҍ^����ٓ���4����y��1.gT1�~�J��
qu(̥�g=Ļ��1[\�4ȁ<r���4�^��1���G��V :�suןmx@d�Yj�7��
d0���u�������E�?^�\�È�*���[��[pm�	8x,���dN'�Vyx��}��i�8�#L�����u�����8Qu�v�����豣�(�A�m��Ia������}�t�ݾ���oqu�pͳ���ie������r�Z� ��~l`r��Z�m:�H��F��.{Ɖ:p]"�k:��P>��R�[�C���<������G9t��pc� FVc!����c�M{�@*��w����pu��Ŏu&��!������S�����8|�KNQ_��1D�@$Y�Q.`�Qmp��P�H�p��IJ��-MP٪C���$x�Nݳ��+��|�vh8��ryul�`�(�$pU���)��`�(&���F������ܩs��+��3��5�U�V,�a�67�
��.I��{��r�?�q�E҄aI�$��s���o��߰��Ω6h*��Fw��������7q�'mJ����o%PN7H�Н�ԙn%��K?�t'��o��rM'���=���|��s9~}�Vs��y�h
N=�PRx6�"|b�@��$$w�C�� ��,�I�A����9�n�v"9�?Z�:Z;�Xy����^�#e���>�l,�l.s���?y�s^���yp��yʀ�b���)[{�|v��M�Y�mN
1:�)�r$�ivr..~z���с���۸�ҝ��2���+�g��d9It���,;��Y�ߖ���+�v��y��v8wG�P��B����;�!;6S���q��[rY+i�V�ڻ|Rl�W���@ɸ��f��%P׹UL �2,>��������������rszZL�Tz��\�̑����d�u�n�lCn%����X�Ȓ�VBi2R�\1@d���uTpX�.�CAf������_�=��n"�om�Cd9��8-�1�ж�f�j�!tdQ��8w���!�)u.�O�+��[Q�.
9��Ӳj9L�7�ަ]T~�Un^�,�w�}�ϕ?���X8h�1(87�pw�\�C1�_�[*gV�Z�	�23q'>$8�������ɟ&������x�]��x^o�SIa���p�.����#]P����b����������nŒ�p�����mY��w0�;��Wy��M��D���I����?��?-W�ވM�n��PH�=��3��1���9�D�]����zH�I}Sh����!�3�X$��g���nq��틤�k�q��� �S�l˙�C7�I���ř�Y43�(���V���P'Q�N}ýu��rzURS�P]�b�"2U�F�7�ˑѣ��k����2�/��"`�+����S	�I���I'��H�h7>��W��t��o]�g����߻�(j���$��
b�����/qGk۫�ݷ�Fzjr*��@>� ���D�rm�����٨�w���Ȧ_��0ߙ^��2�� n�x��������@���Ա3�[�0�����ʑ!�jXG�B��d��|j�*�;&���!W������L'��]�нn��v���9Y>��w��xf�8�gl6F{�˹s��x�<~��r��s�����^��W�"WDQ$��A�l]��
��PE!�ho��{���w��a��q���`�~���p����;��eu� ��=�\��~4I�����WGa����
|*�Hx�7\�껉�꒸}gx�i���3�j^W����}sK��)�엸i���.��Oy��ڳ0֪ܔ��lP �C��N�M�/6Қ���
$���i�y�	J���~������D��W�T�a7��=r����Ѳ:��{���P�ü�~��&�P"d$�W�"�z�I���-c�����9��'k��f	i�z".p���>B~�r��q�Q�NZ:��J�y3gyj~BI� � �W�j_��W�Ӈ�:���w�O��x�|��ϕ+���:��n� ���ݶ*;��Kg��m���5B�8�$\�.��۰ģ�����X'��L�f���X�ż�������{��f����nz$�P�S	��m�#A�!�ފ��C\6��8�Hn��q����U�19�,�i�,D��j�1�?��?���W~�����XH���c9�ti�vq��w%wX{�Z7GE��-OA�Ր��B���å'XY��q^��o$�z-7�|���r���rmu����2���7f�x��N	��8¿r�%T���@��;vŬ�Sm[��E�bI&�Z�Q%D*Vc�l=���_�T^���+�����?U>���R�c���f�GV��Q�����m�"���$��$�H��G���o�mx:����.rɠ����t��:�2w?��J����1�{�=�HA���D�C�×C��3���6"9\x��?�������f�~�q�݌�yq�x˵>�|�	��~����o�	s+�y��������s�|(�^���в'�c�d���	�3�4�Ԡ����v���u��%u��u.�����/��bl
�K���433W�0����r�0��%A�z]rdvv���	U���������gQ��L͔���'������5�E�Cr�3j@ےb��ّ "�hu����K���e<���W�/�x��t�Z��X�	�7�
06;�g�7��͹�scas +CW�)�ݙ����p��;�n�Ww@�p��
_�/�t�A����G7�Э��2�ωc/�xx�z5چ1�3��9��|џ��(q����k�ч���6K����(�����G9�Z�D�6�[foqn���4� ���Q�@u������6�*���B�J����䊇�7��� ��u�2���MN+%����rm�R�m�pV�+P=�+ޑ݈p�h����Ux�����ӣ�f�,3�`1�=�^�/�˭����semv�����~M!��N@�4B'׆���*p��l�)�C3�RȰ|�E�l�SP!R�%�@"����Ы�6�@(�Ǡm&��������{�?��EW'�:;�� n��D���M�ׯ�o�>ӷl/?~�DؖhPW&Y���I�:��]	�^L�q�.�Ѵh�qu�O~�g�@�_��B���rQ��
�����8�����`�:9�8�e�9{r�v�u�v�89���v,�$�5�5;�.���)3��<!�Ц0�BcA��m1-HOi���s���@{�� R������-N�rG�m�^(���*t�k�9���enj��$��K]��n�W_<_Μ8[�������/B����֨1�C2�傰Hx�{w\�?>��ѷ⸎>�>���7Y�����9V��.(�����k1�t��a:[�;����{{�_��F�� ���'��1>�qژ���I���.@��~r[�ɩt�W�~W�.���\�NXݩbz�:1ar�U������+��e�~�B�<�2�|��������=�=�`�eD`�l�GG<{л/����M�£���`Yx��V_�N�k���Ӻr9��tX�EMm�Ё1bূ]�T���U\R��!'/�.����L�Go�o�������3�q�do������<#&���C��,�;i�~�t��&a'1f��~g���δ�[:G�A{lR�Q��3������G��8z1�o���M���#l���Tv�+*�99���M��`)k��h�qXAiu%ʬ�iz;��@|K$	 ��[�t	��9|Y?;�������{��ʅ�O��O��|�|����Ӈ���p��5�U�O_A-ȁ�twޯ��vږX>���[�R�S"���P��z�0����j����xD��Z	Z�n!���'�[�c��hUa�dvy$1slX��D�_�*7�~���w��$6�k}hHʟ���J����[�>f�fѐ�}��}��L+>�	�8�Ig���^�y�����/=v�"�i3ú�    IDAT �U���k�sit�f��E�Nό�7��7q��9*����=0\Ua�"�z�⎎5&[]E 8�����8�k�$��0�m�,���@�5� �@����ջȗ|�5�C ����st8��|=n-'�����_�u������ϣ޷f1�Ef?:v���2�Z�
X�� ��H�؞�N2��٭���v�7��[R����TL��G�:���/Y��%�A!h��c#�GG2k��1�1	��1��0s��ђP�k��8�Z)�_�\�����l�{�'s
:ê�C�[$��wϰ��	�k�a�'�2M����,�g���t��;:*E)�_��,�tҀ�]�5��v�|L�eV�C�l�ݛ��Mܫ�g�8�v@��ɕ�]��z�Jf�k��oSQ7�J�:+nc��6'�9�����o�3�N�z��(2�#��۫���3�~�)綎��^W��k���I�W��g�?Pƹ~�{$��<�h�=�-����5B�\*�=�,�l`qG=)|{�o F$E�Q�_�.T�Zo��h�f�����ǎP�4v�vR��͌-\}��E��l�;m�V���k�[,V=W���s��P��_��r����Ԃ8֗8��z/�]K탸rgRQK�0�w�~�~	_q�8���7��UmȎ�p��0���*T?���e;�vtpqI�J��[{�}���rWo��qnr��~�#)=�Py�W������:�买U q*j�A�' û6V���1,Uߵ��jK�=q�����{*��u�1q]���8�)�1�Xj\^^�ʼ�Q&�p�|�/��q������Q�X
*��'~ۏ��ZъL��dG:mV�RdmU@�#�ڛ��8w�BB��(���3�5*�o%^\[�5�י@�[t�5881bċ���h�	��j�*�`X6�z���Wb���ѳ�y�>���,M"�@��u��4� �0b4���)�#,�Pߞ�&��*��T�Է�ť��N�藿kN���9_�<2���Li���\���ҁ
	����#��#�8���o��M�1���B�@T�B匮 ~�ӟ�=�w���!����R��p��r�^䅿=4�@��	8�@'����N'��|�r��(��	�ᳳ��� �����G~�Gʷ|�{��M�e?ʦ�1�D���̵�r�vc��$�z�v k���F�h�	@]#��#�m5Xyny\�g[i�Wީ��@�|��Z;�Ҙa"�06>`����ȝ�˗����Z�.���W���>,7�7��>^ڳca��.x�Ս�a�a�2B�p�_x��~r�7L���~���S�y&���8�R[��<E��l�oEH�9��]��1�ƚާ��ea�t�o�~��?]}��^����'!}�W| 	��9����V�r �z�(�Z���I�� �hq�S�J��-_������S�
�r�� �E��c�t���Yn��I}������s�S�Ї>T���/��� r�Tg�f��'Cf_Z熭��r��58�������!�@X�ǗW�P�y��u�Um]�(KH+hX�]���u 'J=�x��υ#���jL�jh#��ln�D�k����Y)���	X����K��Ƶ����kat�˽�aC�]�ZtU�:G�g�8z.#r)
�b�ήq"QJx�'����6f�ڜD�针�	�����myvj;^&碘�^�vS����I�,G}w:ӢAi�1�60v��M���n���Y����3����~�޳O�ɾM !"�"���<ATP?}�y~�� *���""��""jD6�����ٓٷ������NuM&<qC|/3V�s��[�N�:u�)�*��@�f̘a x;�Gf^�L1���p��0��*S�*�@)Bj�_=��}2��5�� �@�>��x��pd�����m�s?��O݃�/߇��aG�V[�S�ftӛ�E����d���0٭k{�mm�*ca�����Z-����ڱ]�M�1��W�`[حl�c��k�������]���Q�&!���m�ZI8P��.ߪur_��yb������I�_Ӈ�;�l�k�`m�?IFB�$��aX��i lh�/B\�g��B�p�>}�b����p/��<Nm�lH��Ƞf�H�c�h�g\c�$#��1�X,H}��g����&�S���(ekY*	�aS =F�o���"�}(�^)Z�8�j5r w��ÿ/ @Q�O�eQBCC-�5��&�A��YS'��l����>[�{�J�|��h_w�.v�fN1�f��i���]�ZvS�dqS;�����۰Z���F2'Ys���%�B��T��nR� "�A��t��#:�X�qc�\^����lB�����w˖��e���n�ZQ/fb$x_��̞�p&��$|2�30�g�&ZA}����
ভi��j�жCi���C��7���jy��,^��V`��<`]q3�3c�,# �i8��H�1�Y����Vk���/ܬ��(�SӵЊ�}�Ī�@E���V*��b@ݹVi��7(iQd��M�J�l�J_����>6���K�c0�9
�����>>qƌ�V._��~��t�[Np?�lft2q}�6�DeЏ��aNGsÎlھQ����."�W���+���=����y\)�s?�q��b�䎢��ӭ\�B&`/��L�F���g�*Q�35՘hOL��q{9)~����� SE�o3G��N��6��B;���#<��q^��C<��e�%~צjM
Ħ޲O�n��p�W��
�	�ia�=�Jz"��WHH���H����:/_��-~�b�: 1���P�,篋�s�#����c�$]�Oh0�6��
fqD�U
?��Nު4�5.Ƹb;�N�C��7��l��J�%H�=x=�Cq��ޙu-k_pW}�J�,?s���s���ݼ�{���R9He��)7�]m��ݞs�q[�U��ތxou��8�-p����e�ڠ&t��d<Q�~w��܅��HB|g��8i	�RK䇮v�s1U��9���[�P~>m�P?�����aY�څv`�=��N�I륞�O�����m�R6��4���%nSIgFz�I�`�`��:�5">Iw���� ��:�#�-��	����:�τ�C���/oEKATj�~��x�buS�N5=�F�D�:�dU!���*E�1B�����Ҩ�w$�o���#�.�	i���i2�X�χ�T������^a���+K���MnӺ�n��M��w�[k�Z�0���1����C�/º9��\1-4���II�T#�+�љ�&Θ,=���ս�q߿�F�ZU9��ؠ�E!�~��a�����Zo
�,���.~��扨��6Q=���.�X��-i.J��w�+�!�V�Yh7��M�=�.�!�ɕ>�х�k#��&�MB"̷���я��V<�ʝs�9�U����kj����%*�-��MPs(y��]��'?��?�|��OZGS�őz44��X/���h��o�Q�Vڈ��\�;;�����ۨ֎�v��P1��� `� [��9�Q�c�c�������#���o�{n�*w�'ϳ4k��]����gO��������uR��?g�\7�Q�2 !'�N��ܚֹ���]��ܺe�$�k�� UN��U[�
�&E��-)H���Tn�CŅ_հ�E���H�6�@�Şb�`�ޒD2h�<`����/~�oB�� �;WvP��cI�@t[�R���������l��t"�T�E��ʟI5"�?^�$K���%K0��97�V��QG�.��r9�8��׭J@yp�a���M1��c{�w��i �h�qa�hL�����#�uc���1�/6�0��â')6�<���'bF ��v���s���7�-�~R��*u�C�R�!�s����s��5:����ջ����߹��G��0��(ȵpI��d1�/�v6P��{
�ޒ�(_N� F"����H�Jڂ����q�6UlcE�1%ڏk�p�2��	�½�m�}�INx'\I��̨SFbQe�$ �j�H��N�ظq�o?�s$:y����=�z��e����/��(b7pP�v6;a�V� ����8M��8�]��ֶ���JZ�B�^T��T ��{6#�Ѷ���ѭᘦ,◑�!�_��?�-^3�#�n���#��CHMuX�@�L\�cRN�5�M��5I��I��2i�������X��1u��ݲc}�K��h
���	@2��KV���`p]8�g���"���KPZ=C�+EЫ����(O�*ՀfЇ�c��o�	�38�!��;�b}� ��ə> ~�@�ܧD{�l35#X��0���_<���;���V��^Jrx�2reQ���k��7�p�[���5����W�7vҡ׬_�h��-���/���"���C��l��Vg�ae�o}K�w��vڐ�ЩPn�Wփ�/}�	!4z��5<~�=����A���"�����������,�_���峸�ܧ��Q3`��@E�>���x/<#m~�p����.|x��)���Oؑ�o�?���������^h���ʇx!��h��Ti��$WbS(�9�|��߫�t��o��X�j-�i[D���Ʉ\��p6��N/����ښج�AS�5��w
G��\�B�^﹈�r�* �Q$�Z#3Fu+$�ť-3=�a��X>"L�#��C�gP���~� 2>��wt��<'���yx��t�H�ѱ�m�m�v�#��Joy�7��mra�@�!��^ yr/��o�B\~����|ݩM%BE����:�3�#=�>]��ۛ���Ӱ���< �I<>�r���z�z�Зs�����	�'�n-�y�<)̛����	$(-����pM:2b���2vc��bNb�R���_�����o��ں�8�=����f���_x%|uϚ5˝peU=�]��U��AE��y_܉�KF��p�6��x�w��>(�k�aT�^�A�U|ރ���u���6��H����,��
K�(�u�x��餁�ڋ�X�J��J��r��C�!ߡ�_O���	mae�1V}����O^!.�Ӷ�T�)�[�DV��t����P<{��'�hC�M�P�>y�Ev��ﾯrW\q��1s����[��Ú��[�mU5:��8��r�UϮ];<���tw�;vn}Mm�2F�R�ֹ�J�E#+ڧ�~�F\��fw�A�ʌk����D����)ЎΥp��ꛡ��*t�n�b7C $\���� �͈V����f��"U��a�B��[�6ќ
�Д_�	1�'_iWxy W�����y�锇ϋl����w>! z	��(��6��ƞ�C��w��� ��@эrkVG�4|L���ǋۀ��ߣ��_(���{ 3��4l`)�z��>@����z҉v�rq��s��3 I�XF�)�,z�V,_:�������`j�TxY��c�#7w����6o<��d���h@��߰~�I���U���f���okb2
��0�;�dxC74���}���ǎo��(1����g?�'��C��	�����j��Y�z#�3��"�~�wLLi�l�X�6ګ���P8��0$������h׏��P~�tBk��=��c(�6�x7|H���9�x�
y�+�x��g�P�@��ޡ����Fe$Yz��s���Ez'���/:�K�^�k
��4 N�晪ں<���_������դ���ƍyC[[{�SҢ�9V]���:}��ҧ��.\�����-]���ߦ��v��14J���M���#�^��>�w���\+o�	�ߐ�k�> �D	��sэy)&<;�8Ȧ�_%����-�Y�ٚB)"5b�m``v!?��(8��N2�?(���" ѰbW
�hv�����wf4"��*߭a�o��?�j�3��&m���feo��� ��� ���K���	��v��$/�� �+�o;�dw�g/27��W<�>���j-3(޺�ĮԌ�r⤉9�<���ܴ}{W�x��r�]�m��9��L�tuA� l*͈c�
�u�;����l+dt�YD��^@�ݠ�����M��ڠ
Kk���yp��SR}�,�w̀�:ȏ"+i�;�� ���K��<C�����A�aU���G:�ҳ8�2U�D�	���n�o��)^����!~�P �U��B�֞v�;�	�r�W	����!� ���g(3}����������n�=���Y�����K��!Qv�7�|_��i��v�{3�?^���&%Aa^2�\p[�ZZ�;v�ٽ�}Is��Q�s�H��l��
������>�h�N�u:[PqӒ�$�X@y=�Uq�dƘ�%�Q�0儂��*�k��`q��D���aZGG��#�H ���g"2���sI����u�Z���H�g�a,`l
3Ċ«{����G����TЕ��E9��It/�ɢu֬Y-�@���S�eq�yi�o�)92�"L;����VL��1՟�_�#	��@���o�'芪��D� �pv�ڴ�|m�(���:�Xw�g�w{/��m�l~�Ε5�Ö��C3;�I�#]�H�x����2���ZV^*7�Qinz9�������M.�w�[6o�?4 8ؾ�3�<��pS�Ls�g�v�-RJGY�F�0�v7��~mr0���(_5�"��X���8j��`<3�*O�#��p�ƥ�hX���*��.p�+y� �H�lt��k@!�cpϏ�!m���(��=/Q�0Xi�<��Ƀ4ѫ��8e������w"u���׿����/����g�,�A	��ߡ/�o�N�P���wW�0(=��>��O��|<fc�B?�:�6�����I��)e���s_�Ǚ�g�5kֹ�|����dmg��i 0}���Y3۶�m}$Z�<���QnY��@-֟��wQ��ڪ���2�jV���\�b
\�(ӹ���k)UMp�z�{ӛ�h���Ԡ"4 �)P$�*�N�s�0��������i�Iƞok�H�8hh� �F)mu6�E/
Б�7�k
���xt,���N:��=��i����W�SWD\���AG��l�|�����g+�myNOz�I>�{��&I�{���3'�W�;���#�8�����i_��,}�~xR�A�&� Tږ2��b$��7;���*7m�;>�~�N�p�:����k�ҹ��/o���V14J�=Xm���Ƽ�ql?�|w�UW�~Mn�ܽ}�K_4}����t���1��@[��R����l�䶭��iT1����ǩ�y{�ho�~$R
FGұ�ꗬ2���;l�p��5��O��&O<�[�z�Q�5�AP+ާ����AB�t�8��À ��Q���:���Ω,��-F�w�а�$�ƥ�hd��} @��=y ����8<#�.�	W� �3EB�)�����y�T�Ѓu�ƹ6�_~���ww��wՕW�����HaG�.������|��2�#mP�bEhDl��U���ȍg����>*�=Q�iO>��jm.��p�u�}����B�F�mG?.^�ؔ��򖷺����j���;����W�=��P�G\ۨYA>/3�����ػM>��}�Z�^��~�7>Y�wQ���e������ܨ����\s�Q�{�ױ�y��w��4�c��g�8��FU# $�0�
-vD��������_����V�����PT��0x�@��i:�8af!:�(�ژ�����7H�,������	K�i�{�+&���?:�}�򯻷����_��Wv�4��^{�뮻ζ�i��jX ;���U?�rئb�P��WU|[C��c�%><��M�tc |:�q/u��S^ ˇ#S�;D��>@����裌��r��c�=���/P��V�[���|�?Z=�<^��w��xACQ�b\��\ݘ�/=�賟&�%�����G9.ױue[k[l�dӔ|��( �w�,�Ot��'����u���曭�?աMXg����;42�Y�CP�!:��E5q�|�t⡍���(
��ŉ<���.    IDAT%.�f�G����%Б� �b|A\���'�&�Xo �)_1��3<�Z�����zL�֬Ycu>���ݯ���hqp�s�,H���fР���o� �߁d[�A�E<��C/�6����L�e�.�����ϭdXM�1�#.�ǋ�D����3����=��#������K/�T���;�:���M����f̘ZЦ��� H@����g�Y�mx���;���y���l\�����5+����?���鞆3**�E�C�bR���}���w���E&	�M��j��y���f��F�q��׫$?4�P5�2��K#:�1��s��cu��z	p	������ACU��iO���r>��~�&O�*��lQD���ܪE�2ҭ1^V�D�X,�ʆR�FF���$�����~?+8:��lF�r�n�H�}*�:��a�%e9�$�<�� ����-\�-ƾp�76�\aWT4k/�m�%��LD{QOlߞ���Sqi/��x������\�][����fs�{���I��<���OD�5"$H�&O�T��K>1P�~��[��X֊����_���g��w�x�#���LM,&h4kD5�Q@�l�HTԨ�xB(��;5E��Qg��ޜ�s�w�w���T�$\{��M�qM�4�\�q?]k�V f�� j���#�'Lh���Z�l6��q�[�l-�>{/4C�O<>�tu�
��>����`ĵ:���L�6�\�M�6������%PM�mJ<�Q}�<� �Clk�|ł,���3%PV�V�
%fF"��hW�E���;��$?���ޡ��*N��{��xCפM]!R�3V����np��w�6�5�0H�������96�͛z�ڵ+���/˩׍�I��7i���p�5kW�|��m[#P_�Fcuε,}n@�i ��:���c�ns�Q�.�H,���J�ƯQ����6N$CEC1��kz�, ��x{G��� �iej����R���!��)�t�kש���S��� �Z�\��2`��z�Ϊ5f&" �C�K.�� �*��cI�Ԉ�59�(,�j�~®�&�ŀ�|�Ȱ�2��r�f�@)yT�F	��D���
�;@*vN�!��A͕$�`��q��<a��C�@�tY$C�#��6����GlL�XCm֌K\T[�',W�C��3r�F�-&L���k ��|O�s---���Ǘn؍��cO8���r�-�t(���sPǤ��8��JkQ'������� �dƵt�)��yh7Q�1Ѡ�5k�{�ey�,�'Z��qXV�#�b
%�D:Kj��%�R�S�]���̵�~a�:��r��J���+��j���n��vsO=�4��u˟]a�b���SO��ɛr�'�ʠ�J���nӛ��P07��lJss�V� ���
�ZIn �� p��ʀ���{�����a п��A/W,ā-�}ڇVD�mV.7D%���&�.�\���u�N���ļ�(`O�P(�т=c�@�ȗ��]�:���׃�����'�t��h��x:z��GVJ�U#���8�U���o:��LWϵ�._��~Z��8�"0m4m���\:�Dj�:ₕ3���l�dĚ&Ŷ0ʹ���$���h8:
j�t �y\���n�k=`�uWf�h�C\)�ػ(��1u��P���E����$�$�㘖0�=2T��Fٵ�I��5p�� 5�A@]&��`�g��α�خ��j{����[�� k � ��R��g����͂�z���\J�.����Y�ԋ��} +�I޴ruf�4����f��n�?����c�-�F\ڂ6�p�M�HV�vƫj�(��)t^K9D <I�����b-^��I�
.��y�-Ʊ�2%"DW�$ �`�k��!��Ih�چZ5.�����Phס�]�N$$HS�?jx:DJ[� 
�#�M��E�i�0�����Y�� �5���=�z�f���%��QD���1t�����D`�v0��pHhc��N�(-j�Y�1Px��X��Y7u�4��_�r�/���0��Ǝ������'?$K�I�݊O }�J~�5�-��5����@�FLh�l��%T��}Zp��}�8e�;��jfEzB��5��wҧM
��7�[j�0n�
{��~��6�_��K�ɿ�׶
돯Y��
]%	Ih�����y�鿘�J^�e���p��]j�Ff;������-��M�Ċ�)M�I��]�Ѣ�]6��Fי3�A�ӭ6�.��$^b�t��Ӡ�^	�`���(W���s�6�$�|�E(ZlZR���t ¢�GBj;�:
'�E���O��۸р#`B��� ���>q�JLG!�G�.5�p�#�p9Q^[�T�5Do��c�2XX? 0@�����= N�JE��0����g��ͱn�]���� ��/�-b�4mH{�1��o�f��d�(��k3"$^[l(y23M�>]�GcV��`�x�DM��K����.BQZ�\�(�\`�Fe���W.lٲ�$�R�������U3�l�u]}cT.jeRTZ�Z��h|,3�F��(T������RZ(�t��`�|&L��R���~���M���0=�e�K' ��h %+13�@u7]nu >N�i �CN?�t���-}(8~����<�V$��g���"��Pb_W��C�7�����كrM<�H��1 "6�o��)/�@�'�$ġ����� ���m���6Ȉ��A��[�Eۥ�W3'�����:��9N�1�͊��C���ؠR��I�5U�d,O��w<3n���כ�E^rׯ_���/)BY%��?�����mk�����\���k�xݢlw�ɢ��Ӷ�nk��a�ZnLݦ#.P�ǃ���c-T������f6Ow۶n����H�; ~Ş:m@i�((� ���\s�,�`��MA�+I3�Du�J �)Q�7J�g/�"�N�P���QZ �a_��݄qM���4��*�7ʁO�dJR�'�ڀ�A��ZL�2Q�4KH
���n����OSovq I�R_��.�jm�igX!�)j�3��0��8$���?���)������(�~�d�^���꡶�k�'�� �L̫�]/�R��J�T�֦�\B'B�$��=.���P��+�z�K�m�a̸�wvl+��O��{dk����������G�����/U���Lx��5���>h�W�K�To�^%��Ɓlv�<�j�.�%a�ĩP-�Z{ń:�[G�3�|���[Sʗ�s���/��\�Z�����h���AuZ..W�%]'d����fT�xA6g�~�m@�Դ
�:ƪ���_x��c�ug�u���<��%�?�$��{���c���QQ9ׁ�񌝼s�=�(ã�:�x}�>��Ύ�ݨ�҈׮]�.=�B��H�H�2�~JN�I�����%�a�A�U�1��)�CY3�|����O�W댬6��4 -�V�*����KZӈC�����O�j�:Y�¯�b�T�Wi]���:�oK�}<�7�5�*�>>ߨ��m��=���6+�+���r���m'�,�硕�χ�C�L;h�\�O�+���@�&��9V����+n��K�I�7Zn��`���c�ĢX�L)��EK���.����Tj��9�>����\����D�8քGb��3�ȵ��VJhƃB}YC]�ĐMn�n�ݶ�[���𗀊 8���y�Fu�>ޣx�4<.W�z�ᇭ<�8s�̱��,����B~�E��A�ZҜ�҂]+Td���f$�-7k��K�s���<:�����{�ԋ���Tߓh}��y�0�K�j���r�C�B�p#wYn�>QP�JKg��t�l\9V+�A~1R����v$uPO_n�]��A�#MK�������ܟJ[�=��)�
��w�t�#��Y`a�klH�/��/!/����&���*^{�wݛ��&��J��U0�2l ����;�t�ˇK�X ��qPK�  �C�����Pe�b@��98�%-���w<Pn�!Ϯ�7s�L���'#
e��9�`]����wG[:wĦ��Y,Ԓ%:hs� >��I�Q�yqsjr�y衍A��ǻ@���!�r�O s�����r���sҢ�ob݌-����X�G^�*,� h
�?|� 
�x�� 4���$M8(nN��=t)`# -�yo�	%��yy%~�|)�>�校�(Q(aӦ-�����'� �tI����*)Me��e@��������6Z��i?+Qf$�NKڗ)$"��w�+.���۟��%-ٖ���x;�m�s��Qn���/>!�%�}ƿt:�2c@�=�U7^W<8��AS=@%.�?,(	��|� ���Y�_�$] Gz��u&�!�ǳ���fj�s��@�.3T���hv@2q�%���@�I��!�!Mޡ���J���^�k�i��6R�F!��64��+
6 �u�@��o:�3@`�=PE�lPN(;ׄ�|���i���
p�C������ȼ�=*�lİ���,bаI��t�g�P$�:3^"RN!�Ʒ���N���/I#+"���X^P� hX$@Pz��H�C�uHC������"V���g��E^��ͥ�3��f�pq
� 0A��߀�Ai��F�u�*�;���b�� =q()�!�]���� ��&�O�
� ~�(6~���9Zw�"��-x�C����^��8����klG��B9;ޡ.��@�2V��^Ң����;#�Ϩw,�#q`�Q`QUTI� ⷝգM`3�>�N���`����߻Uk�s+�[54` -T�h�u�Mۼ	@n�YX�[�~;*����\!'~^�4X�p<��g�5!,P�@+�u������}�r�!n�=�k �8`�ts]+�p��Q%���pV�6i�^�-X��~�h_t@[ݩĎ����1*������`�s{�၏n۩(��FY+�o(���u���(p7�t�Xw̴P���Dx�B��� eo�%&]@�~�9���f�(��HCڥ��L���,ΦM�LJ��%�}X �֬^m�ed`Rn�3� �*�;�Ϟ�d��P�4����iaT��gkOt�����m�1$� &	�u��Z����2")�W�Φ�C�k!��֦�	�tmã=��
Y9���Gn,����{�<w���{�9;��qh+F�ZB��cD�v��}�_@��NgD���~kQֹ���H	y�d��j����;���[�l�kٸ� �gH�P�B�	G���ni���a \��k���$�KV��i��>�ܭ�-[�g�>*����%��$PK(��ν z
�̢�{H0��h����=��Z75���1��@(��G?�Qw�܅a�x�7Ņ�By1��;�-*��72;�Y��ʿ���u�]v�{X�6꿇�v�ʐ�2</���}֝w�y�e㝔t�}�)�g����neb��AO\��&��䟐q��wΰ��W��^'�C좶�D�@� > ���������Pn��vQd,�;�F�ަ�[���S����n��V-l[��>�Ԩ���M�ɂ�O2�3(�V���� ��<��Z8_җ:��w�˽��T$��,�Gy�X�F�N�6��m�̰!��O@�O �(�z��S�l*���_�~��IF�Hν�-/��Z�����X����"+�&��� �@Q�Q������Z���}��ƣ�����������S+�'d�7�|����0^�c� WI�Vj��e�Q�a#����tg�}��C<��O>���'-(qBJV�r2U��A��y��J !���X��Td)<E˺3�¨���Z}+JB�����c�] � ��7��K��Ve���;~�K�z�7����b���� �w���<*]f�@D4����5�c3Ė`�N>�++�ɀ���+\ˆ�n�[�w������T�N>���Ԅ{��%Y��gZ�SPo$.Vv�D���AU8�W��Zf���~��!�Q�Nb/�� �`TjK��'��ԓ �o�ov.�7(��-���7��	��	X���7c��in��*v*PR����S�-X�������T��z��bl�u\���3��ܺi�啒,��.W������vȓ�*�f�D��U�F$��Rht���Xr�ع5�N#���2�
���
� �5$>fVӧO����O�4��h��g�c�]G]���OD��%�#M('�� ��a0 Ρ.���0{�"��Sة<���߈zϘ1��J� 4���4y5]>�'��*���5����	�QG���{-HΈG55ː��+`z&�3`$ 5X$$ ��1�eцd���V����~B���S�.8�A'�4	l��f@��d��>��u�ʚ�ubs�u�6�c�9h��e0���E$�~Hh`oX� ?��=���Qg~�ڇ"�(:������i����r^��m8bDՏpaԁ�>�6�[�i�����t: T�5Ā6  ���o>�\9�����($�2*w���b��b�
wđ��H*��(�=���6��#�x�M��}���~��9�����_k[��v��@o ,���x���Pf��~
;���u�;��J�(���'�RuM}�������ʡ�?���x��m� l�`ј���1�@(�"���$`���|c'���*�'��B����jݺ{�<ȏ��/� ���s�.鍗�W�0?'�Ri]r�����	�,��gH[ZZ�y}�k
�>�t)y����y����/KUM��m��,�)���/�(`�Σ�rwvV�(�RbCl�� �e( ��%�;�),
��/��t�����X��J\��Ip�;���C�q�'V��=�N���/����(�9�Am�sf�u�������#�W"��_�t�׸f�(˖=���t�^R���aK&�V��Ϣ�:�3���6�uyf��5
���E�=v��˥74s� XP9~�0�
`��A�s3��L@��eҤj;7���i �@����s��c�I��֜��!�m}��GO�.%i�P/}�Q�#L�1l]{{���?~�>������a��Y�e ��S&ҁ-!P&� [FK+�	�X1q3�L�.�Q6yaDV�/u�6X��f����=z�N4�f �N4����Pp�s_.(��2 ���eQ���ü�։bZ�:h���3r�\%]���z�׼�xnxr �T~Pc|Pm��,qJ��:�Y�ʋ�"���&�-�T6xd��A'cK� Y���C��_�.���喊8��/�mR��SH?�t�Z\D��V�]�ϨdK�2M�ɲe)&����� jz�h�� 0P��ҷ���ϻ׽n�4��
hC�wP\dɲc�)؀{��'Lvλ�G�򁠴��K�kP0S �A:�T�=J�����Yљg���~�;�)'�b��%]�9(�^��w�*y�7����c��)�H����cN��w����-�@-`se2L�PPm��xx�š�o~�ݱr������&��n�M��0 )���CZhb�3F^� dM����W�#`'z��m��D{08�9�S��4i"�����/���c@���H��9����s:VDe����RJ3�����2V�]�ψ��K�MK��,&[�7@`�
���4x]��a? $ �j����S!��}�C2 h��y~`�S�'�m�3 ��<�YCy�� $�	�}�zSV*����a]/y�>	�G:@��;Pmf ����6sDc5X9�0��:�Npo�8 �U�j	��8�{6�Q��\�o��I2e!S�u�go_�͚���r�B��u�P <��q)���R�*H�����v���%����Lx�U�ͻ��|x7H�"�6�b/��_�FMM�ޑ>yF���w�.C����NU���l�ǔ��~ݳ'HM�h%���۫�����r�Hz�G���]?�Np���x����Aq�� �3(0ψ僢c��Vrf�ƍ7���GR�1�L�8��v�H    IDAT7&����2�y?܃�����M����rK�5�<8r�@|�!>� �0;q����r9�}J�z�2BGL�#�:uE"�f�yM���G���I@����6 ��68#�����s|�q���k�I=��qFώa�<�b�]꨸H�(���f��A�M��a-���,�`�`C�Kc� �8��8���e�.��������+g�x�n��[�'+w_^o���W�eg�W�Gz�����d�b1��
-�1 �J��D���()��f�
E�
��{(*T��p> ��/����_l�S�õ�܌��5���\4���т�5z!Pk�4R�((�ɡ��r'L���}��
#�:�����S��V=gqƌmP���ޑ&3��|����v"�Ê
�C�������R.7�dݣܲJ,˩���� ��e��6`� �z�g�����u����v�m�P_n�N��a֬Yn��*��N�6�އ�ت�K0��+�ѧ��W�����s���������t!�� ���Q,�?�Ye�����#�}��,ű��@}�:��� �M07åڈ	����/��L����{�]Jz0
� %�(.0A=s�����~�=����C�����9�'.�q�i��3|���gq�mc|�
s��g�T�0�
�xoX��UU㪙CM[M����}{����;קܜ2�bi��s*U���ŧ�d����R�	��i�1r��F%�[[ӹ�s"��4�8�� `�f���Y�@�=��.;}ޱ�b,
j��i������m� �
o�Q����o~�'Mo�aM���U�V�ռ�sd��*^�ޥ��L�ރ�6m�`,�\!�V��B���ꡛ���r�3��h&��{� ���Jp�K��qݸK(AY����d|�AE���H������v~����ͻ8MFz��I"h�Э^��s�a;�l�N �,6?���L�ì �vX|:�ޤ�D9ɏ2�`�r��x�y@M��C�>�F��O��Jԯ�%R�K92Z*5F����r�?��Rp7'$��PƅS5�  P@��*I?X����:=���E��ɍ�r��!��/��s�央���������Zy[z�j��轐'�JLF�-�>��������7q����ex��V-�\�6r�f@ןH!& r)��M���F)�kd�U,��IPP��/����a�sB0�7��?���N�c�9w��S�����:m��#���~^Rxf��'P߆����|�m��T�����A~�,|'�� )UyP{@��4Zo�p~D�lJq%�)��6�T$Y����m���.F�H��{��M�:g����7j����+iȾRȨ(S	 ���&��5�^owK]�v�}w;�]���i�C��y���FM:% �3j�E�
�<H<�J��$����}>�v	�kn�s(���9���=�k嵯�&�m�( M\Ր%ff�x�H<�L��u�bq[���I��W?�w�
�E��J��H<p��;(�Oj�}>��zx�׭[�+y6σL��X` ��	��7���N'ع�0i�'����^�V_� j�q?�P����q�v�[[��Ӊb��,rB��u��%֡"�L�~���6ʆ�I`ة$����x��'��?�+��`7ؒ�?�e;>�+��b����WG�J06P�z� AG�A�uO���Y�Qhv&���;�p�u�>�Ry_�e�&�enN)�Ydq�4@"^����G#����%����n;(=~�V H�X��
~���.���,��?�pw�G�3G���@X���}�{F�;��tD��')iB]aCB� ���oE��}���n��`�1�� z�D�U�7-���B\���s�Fp�_�$��E��~�'�C ��W|���zM�<���o�E���/��G����*9��=�AP�[����tn�5�Ɗ��F�mSm�i��-J��h	b1�9������Sx�.�f�x6U(i�ғ< ��N�1ʾc�}�<ŚT�pCg��0J�Mח�=��A0 x0���;��,��PrO����p-�Z$*nWW���y�<Ɔh���Ve�8�4��X
xl���q�Ȳ� "��T;���zXy���ܿ��H½�W�34�dJ�Hm!y�8�=�o���Q	�f�+E��82T��j��"
��=؁�@ƂL���5Y��g���K+vZ�� v�O����=�K�`����t���Eb<Qc:)X���X�{ޝM�I0�'"�D�W� �HL������Z�+Gj�_A��'©�F��#�gsz��� �`[B���=)br���b�|��^�nk�]�O�X�}u䳎���P�^�"H%��P�`^���l����@�Ȱ9��=�y���?���o���x�)>a����w�ml�� �� b&``J�)��.�=��{�w@�E��h�fMW�YY�4�t��	���C�<n|���!�KN@�(� ��7΂�="¨��S�dl�1!bE�5����٧"������ )"�^D|�z�:�æK��6�Z�;񤷺3���|N�n�4�d���o~�D�u0*���|b:�<�ʒ�)��+j����J�`	� 1�������à�:�rhu�7��B���0��ފ)�Q��_��Q�!��"�����������P3> �Xr� u|��_�>���X���E���_��TR�/_�V˘ �$�{��d%���x?Ҥ� �|��� ڂ������|���皼�;!@�0�`��w����vC���{SC8�ܥ�2�¨�@!33W���C3� 0P^
�*�>5 �x��ܹ.)����o��g�=c:�����g���ȇݏ~|��#uڪ?P��˔DR���PZ4�2b/����-�m�`z�a�߸�t�!*;�2]�B����}��K�}��p_>����+w1x 8u" l��:��1�KxR�)�}��C~�U�/UG�=���� ���xh�y��^�O"A�"/��� ���k�UW]���PMT[���<p�ZFܬY�L.���,^����	u�U�;q�̙c�O��)����ɓ����a�\F�N^,|��./�(X���{���~� .��R����b21aTR�͛'絃#��-Q����Ȝa�+np �E$�ڜE)��2��x\��)İ=:� �� �/��U��I��@ ��cG��QXʄ/p�_M^�Cz�U���=�'��)7i�<���\PtS�1��|�,��#(�JpK�[�+���K4� � 
((�� ��@�~�[�j`�3{�[��<;�:PȦqM:�}��6`�o&�ːg 6y�>��;z�\y�<-l��j�b�\�QV�y���_kG?i	�����=$@�E��wKd�3ْ�47�y|�ˀ�e -W@��X �"9�+T�@@	P8e���W���u������Z��w�o�p�Q턬o��#�6?)X� #��a 1{�7���<�<#j ���ǥ�W�
F�L�B��d4���%�F�>�T�V�6}�s��@���G#�#]Cq�I	v��� "�w4��2�����׿6�>�ܪ�N_������7$1��h6i�dY�<����y�C���E�Т8�o,yB���A���P77�4�5Y_^�u��R��V�j��0X(�^r��3�$F�#崄&m0R#'�Bpۙ���NG@9��w��QP���b\���\Š�nYڰ#�+m?΢D{�Z֭qW\q�m� ��%Y\'�~�NF����h@�� -�bO)��	f��k�� ��9���(�ǈx���l��MF�I�4JJ�r30@U��@�5�C�7�U��s���ߡ�sT2~
	w��(�RM����L�4��f�mSE @M0Ê �`�P��8�?����7�k|�X �����J ���%�m $o�-G(9��������{�x�bs��q�y��,���~�ӟ�Ye�]�~J,3ԝ5 y��Wyi�J�U��
�#:Hؐ�J�e���_G����Sj�����&H��\A�?� ��ȗqd��!�e��@�
?�;T����F͗�� �8q�Qq�p����G�1!c�$b<��y�)wU�9�dNI���7h��j7t�[��1�-�}{�vw����.���::P�4X��؏��zP9�W�A�_����x*�M��۴|^)�Īd��吐�aR�^��BJ�������}9���\9�e� 0��Q9��v��x�8�u�򖷘��I'��6h�/��3��#Pl�Ǖĕ���	Py����;�^z������w���E���Or�i刉�&M0��>8��#7�%6��а+�	&��E3p��7�{D ���EF]hv�ڏ�09��K�s$~X�q?���<<n��`SPl���(J?V�6Y-,�daw��xPu�3hx�4����M�[B|���̮_ߢA�^JW�R��"����o���9��Ӄ�׃��d��z���H����ϖ"^ڮ4�X���0*)���zmF�n�'P��n v"�y�t���dܘF����N�����Κ5��	�2(ؕ������%�Okq�H㩧�rϯi�"u��ڨ��.�E^�<��r�)�u�}��ݯp���o��Zm��R��+/� '��R�4pٝ�+��r]]>&Ǵ#&�Jpo�V�O�Q�K$������\Tږ�ڂemW���=x�*�'ݑ�ι����^�׆/�M��dQ�}L�@Vi j����Vz���㮷+�>t���S�~�uw��"�3�p�v�����m0��e�0�`]�'�v���)�LJ�Ȭ��J0Lf��o*�ŒD�N��L�$)ݪ��8�]Y�d�;۶��0���ޠ(UL�~��9�sg�)½��p�2˨�Ă�%���;+`��B��x���ũ�K��&����������"�=������xu%-L��ȏ`���Ǐo���	�M|t��|� ����@�=��<�m�l���D��g�zxgW��:pO���FS/r�L�\('d���et:�ۀ * A�l�e=,�@��K��K��J��q�������e�N##����7�!��k\���ɛ���뤴-[����֚4�<���Nw�]w�^#�9����{��$#c��z��d��l��tv�[�h3Z}�~zqG��]�-�-K�5RNE��VI�c$�u��j��t�$�G�O����nE�fW��Nω�'ϡ���PIuȦs:����KX��caZQ����[����T�k_����"TT�LZ��s�����]w�Ҩ9���
l��j1�f���t%���:[�º���ڀY	�f*���/�"ۚ�4�s������ۋ���Q�͛�����������w^d� Q��. ����η�==�A*�A0)|����NV\rl�?0��@��ء��ץj���Z9�!-Ψ���eu�:x���f�2��4F�6	����D����?��ΙG�����@�Im�)b�$�����c~�F���D��=<��>���_�!Kl�$ئ�Uq���!�30��p�d yH�g|X�A�y���{��ܩ�u��`(����	�	��
�>����<�#��Y޴�o"�M�6����m�c���G|h�6�[Le�]��#�x�nxpcY�P^�[rv-j��6�["I� Y~K�""�ۨ�vu͉L��>��}�1ڃR��Ϝƫǡݺ#��搠Lw���5�����;44��^���y9���{��,��ig2#�Tݫ�j��(� ������wާM��6��?�cF��]9���MD���0�LŢU#���$Sq��)=�*��g�J�#GDƐTTŉ�b��v�MV�K��(g�>۝��[�]�����.[�����i�2�S`{����C�PZtLP�x���M(e�v+�;�=���7i�4��B�o��;��xagV^{ݺu�!��a�抂�1N�	�(�d�	�����E?��6w�7ۂ�����9e#UB��oA[�|]*�j�N���xD6Ŧ���N<1a��[��u��~�S*�� `����d�P���^�	���<+��E�<���lP��:�v�W�8���;��Gf+��W�O\��u�Yn��yn����c�u��DVi��U�쫁ǢW�M�x�I"|8�P�/�%1�C�Ć����L��zW��fiE��m�\i��|�N
���(w��<E��Ɂ*0�7����$��_��W����A�9��j��vj7�{�ᇛ�5���܁j���<x؆g�%��'�x����Ysܷ��-W%������� �o��-���ƫ��=[�9�����,1Pq��D��P}ṙ��8o�������u�܈�RG���e%�<a�ڶ�� ��v05�3�s`>����k��.�:��G��jɣ���'�x�]{�5bn5pV���.�HMM���Y N���I�y��2��<��3,�s˴-��C��"6�*�|-n�<Xi���8��*�f�2@p���1�侴K�i�%C�t@N_��F�#(�R�-y�h��W �ȕ ���9�4��z$� <+���v4��O��S�)'�͜���u����`��G�Zs�5� ����<��'+��bTP"�a��ꫯv|�!�5ig����@e�kN
V���J��d%�ā'Ѫ"j�?�!pbH�Sn�x�3b[�v4J���^G+��+)Z��I}D�<����N-����4�ۛ��f��Y\�yƙ����=��f���}��Da�lX
���HW��J��Gu�Q^�5�9�2���v���)�O�	��W��v��6v��d�<�/��^�,�a�FL����hR��u N4�Hź�������V��W%%Q�,����kT�6 �Tn�2�Y8r~#@`��z�9�8�(�;�\���w�{F�0u�]c�V�7�1�q����x�������w�_~����Ns�Y⹱��w�}L�kì�A�ƍkl	�ܤ��C :��UZ߅cK��3D�1��r��n�=/?�����QJ���'WN�X�BE��y���C���hz�+;��$��5����-�P�u�ofc˜3�<˵i�v�Drx��EÕW~��a����Xޠ�A�Ix�e��o��s�=��ħN���XHH���{6�J��dU���p�qΖ��ճ[�bMT�WR��f��^�u�Bk���.l�?*���ԇ��_�JW�uؠcz�:C�q��w��3�">��;�x3F8��%^�Y�R�&H3n��FY7�"��gFJ���/h \�^��W�Q	��Γ�p�6c ���R���g?��QO�)3;�������L�H4VҰ��P�}�`C��ŋG�٣��'�ږf�̍ʻd��L��Udق���E@F/C=��%�@�˲�߼������|���w ��&
�����E�v�Ĺ�R��㠫MhsG�'�X�5ԍuw�u���W�po��7��u���Z�x�gW>o3I��(�m7�%�ں��xB�`�s��|��L���z�r���_�E�#5�4���-#�x2'&�ɘt�����a��w�n{��A�*����΁B� ��� '.l���z�灳}.�Bг1�]��l�d�yg{�(��� �/���'L�5O�΀op7�p���n�r̙;�]t�E��s�������u�v�$۲f�x�:�ր^��(#�0ȏ@���2����l�U�Tã���������Bp�ism6VG#%����~��%�\:<#�a���W�� V� ����>QO�shp0H�o٪���J���?c�N;�Ĕ���Ci�0����f\�����=���n�����`N6�o�$&}n}�����g\�FR��2��'aP�'n(๽��zl�ʈxH�ע�T,ǤӞ��)h,�\�Ī:"��Jp�ߝ�����RI6�t<����7T �lap A� |�J�X    IDAT �/}�E'*<�j��=)�W(:���\���fhx�4��[��^{.p˞~Z��:���%��K�R��W �.�T�^����?������(0�G�K]mM���V~"�=e'��C��pWWWe�\H�k0ީr$�.E�Z���0*��hM��3#=�m�<�έ:�`S���7�̀�ā�#��ꐤ��z�H�Հ�+^NԳ��^[��A�⮮ќ����	���wP}0-TEȉ�K�ɀι;�h
�� Z@�����m
E��n�f
U�����m�P>��ͯ8N2m�SbK��k��:��}��k�L�+j�s��;*���m�O(����JP��g Sw�uD��,9r��[l}�]W�t2����>W|r�d��i&������Q�-
���#}@K�Ȫ`�Ƣ��SNr���g�#߶�E:.���Rռ��K���X��6Uq Ȥ̼B �ؗ*�Q�蠺c\�)�e#K�W�����,�4�^��
   �^��%�Q]Se�.`d L���}r�v��߶�X�#�C?��9vO�����e��R[�C�D���G^�>��=���s>��&�����%`w�w)mY���� O�:ո��$�e�-Ly[��5�$�_T^�JD�P�H�":f���F|d�Q	�������6)^!���PR� �
`r��*,2m�Љ��Vt{�O����
d?D*�F�Y��@O�֘� j�}[�=K	�d��mh�f���w��5E�{{���~v�]�*�(=R��.��7���}�B��a}!㉼�#����#bxa\G%�{z&�Jݫ�>�{D�j�
*ᯁ���5K	8�?���G�O����x�ݴxh�1t�C�O��7*�����d��b]�.��꼤8�d�_����ϓ�b�5߹�=�j� ��X\�/WJ�-�0*�I�0",��"~�"wm�5�lQ�[�dA��m���(G;Ӊ�u���}�T�o��v(�R�P�p`9�~� *�(|�:E�a{[ �k��n��y�,�p�H�{����j�|挙���	b/Z��&���m؊���\}B�B��p���p�������D	x��x���|��|B�,!�Q=�aB�5�X��∣ޣpA�"=�MD�R�X!&�-E��|�H��NQ�:p	��[�n�֢��f���p|�BXW�~�Zyb�W�d�;O
O3f4�$�o���U^F`dA*��z˛�e��#�&Y����6�p� �f�� ����)/��<5�`--�k��-+�m�����@���h�>emK��bI#�n�b<k��#��\���Wv�0
�]WΥDBc�y���$l�- 0@���?��Sm ��T�������1�EC��矅$O��8�v�-[ni� ��/`��-�k�j**�Gy��K��a�`��=��?,���~�Iw�]w��+N:�t��ծ�u���M���zK�هن4�5�����Ŵ�#ENX@�DҒr$�b���ҕ]ݣ�Kd��G�X|ugGgj	�� ,�l DA�)�HV��
���>c��'���������vy>�� Jb:���(�?	�CI�?雯o�������ڵ����vBZB3˥_��ť��o��M��\x�%��/\�A5Fik!��a`�IT�Z�q�0X����$�B��T90��{�0B���NTNVf���>��PQe� P�+!HF  2n���=V�
h�����i�l�/7MM����x���S�E&�,,�5H�ee�9���PU!�Hl�ڵkm�g@b�U+WH��j�Y���!^��l0�����M�J�����BiC�	<��i��{<�'$��+�r<�!���t��0*�].W����
���`���H ����
O�>7� �W[#����Ǐ�`��p�;��8��)�`Q3V������ g�˳ �h����cB7E����N�'�|ܽ�q�ۦ�(OR�,o`�pȃyT�AI��N �a��@ⷼ^u�;�P^�dI����6��=ɷQD�I�SH=T:�Ѐ� � �~�1`Y����D���^w��6e�[�f�tLnv���&��B���vx��`@v��C8w� ������9*��:���w����̠�XD���y��?ވ��	�)+�����������%�Ή
Ҙ�೬�93����	��r밺��i�bNC���R��xa|{���7c�$���Iz��9�Z\WG����ϚYF	_��W�;O}�9��?�,�$B���\^��;�z�������C�VEnDO��I>>k��֥H�X�-���5JLR�Vq���W)�qQ�I	�A�`����w3�f6"����LjG*��D^*�LJ��u�{ڴ���֧�W�Q(t�;���HI��~��3�k'ˁ�M7�d�ϐK��+_��[�j�m�j�'�S���抁S�8<�c���X�����Ͽ�����c�<�#��VF�LZܣ��7l����!����q�/.��u�Yc������5aԁ;��Z(�38�7F�5⇽~���NlE�:�~��6/j�V �wJ[�Ȥ��Dj�6�� ؂��OMZ�nI�PxB�;��ʎ)]�]��>V'������Z�v�`�}� x���� c� �0H������d�5�M�T���rz�܈�Ĉ�H �K]L[0����1��oѱ��eB��O�^� 8��$ ����d�	���X�[�#�wJ:��GG<�@�B�|�_�e�=���҇gl���I�SO-s��|�r�����WK|�x(JawI��@�\ ^�8~0���&�^��������.��bm�0�G�lD�V��;"P���,��5]��9\tq^,Q54�B����0��zV�<Z_�M��X�3�M&-9�E�/}�2R@>i�d�+��pw�_0�w�j�������;L�5�HR���R�ɓ��N'�9��a��PZ_�hZ�����˟��[����U� = �+�D���*hs>���W3e��R_]}�vF����Ė/_.n�(��v*tDr+n��	���v�g����S�W�F'�Ǝ�wR����y�m)��,������2�3�=��$b59���O/�0<<_u�{z��ģԛ�r��Xr�d2�)[� �$����P�ԒE\WW�{����<q�D㛡� �<�Pf�#�8��}�<� P������X�2��T��n�͞1h(#�D�-�}��J���#Ik��Kdzr�����R>Z[;��;[մ������n�xi�-X�t!� �S����K�5p���/��%��д�iӦUikmm���j���:M��������;���H}~���'F��I��hYs}1��b��Fr��&[j΢�1�.h�!Y(E�3��HT��ڷ%J�h��ݚ�d��մ;�ر}��Ha�<`6�S����렣�u�ف���G:�mj'�@��g �k�q�s�"Ӡ�o �I( �Xe�����^:"8�� .��	����4Pa,�E9�/$ZdJc�|�0��ߋ�x�K���.�ރ-	&�s.����	0/XZ�+�����-ֵ�u,�0cƪ��{L�Z*56��*�&L㸆��]9�ɕF�b,���)�E92k�>:�-�(F��h)Z,um��j!6_��do)2�M工]��N������L��4���6�reK����Q��K��������6�4�Iɪ�"��I�a�H�8�*)X.�uu�|Ok�:^��R�ڀ蕓�Bv SǙ.�BNjrZ�E�E�S�G2����ܪζ���J�\���6։���H����	�C����/O 0 pf(F�� ����I��28|��OVD�H. ,:( 0�R���-Gq��2Q��T}܄q2W�Ii%���Y�:yse���%�	�b�.y00��.�s��M�ԋ:�qݫiH�^�d�ɾ��f�ŞX"9X��z'�tQ���II��"A1���"b�
b��IR��~����b��:]9����<����3��L��*_̯�<����n���C��j�ͷ�?�����/�u���x������T$�O_w�Q�xdL��;�l\?`�%۵V:�¢���v��&W}���޾�v��<�eiF([H൰�&�^��b�!�l?ƻ6`֬��^���
c%,@a�����H�:Ǜ�������5#�[����*�:�ԩS�NUQ<�2���f�8@=tY�G�ճ{6�@2X�fx!�3&K��1 ��wٝ�^9�L,ɨ,Ϙ��y���`Io��r�<��\���j0�i�l%�A�,��d�Rn�����~�G�׽������%=V��l�rC��(e����?x0s�ո���W2����5�!������O��W�n�<�Kc^�W��ԳJ�����ҧ�N���{�{gwe}ue���{�ޓ�޹ra�����k�o��{���ǟ���o{�;~$�~L�����>�03������W�f�F^�v��3�7�����Np0�D�Yx�T�B4��R���	�m�S�N�2�A�uu c�g:S�;�B!�⊩�ػKj/m�݃��	�k�W����a ɿ�7�F6�����S�xO�L\�O׶��]_����.K���ͧ��{�~������o��L��#a��sr���A��{��*����Gԉ���Gg�����EX L�YyF,�����ԭr�����l|�<��U�C��O��4rG|7��Çv33|aucm�����pbym�On���>�zv����?x��Gn��ޓ�W&������<���x+S�^�g~���W>g�Z�gs������qi����s)z7�{�H�Ă�xn6�n�,�c(̍��`!d�"���U�3��/��o��L�
D��`ZK�)&3����~��"!w�E���΍	�$���������ۓF������w��\V=��X]XW�g=�Y�O��O���7}�7��Q�q�1L���!�<]�gTou.���ׯ�i���3�z�6�h1�����i�>����s�v���<G�-�w��jYc�{n]4�����3S�ֶ7ߟ�y��������Cǟ��C�����2���DV��Hq�K�No}Fv�y���Sw�̎��DR/L7�/��D�/&��:�b6�~�U+�a����ǃ��Pq���O�;�R��.�e��N�C��75૿���Lw<'��*���E��QgP��7|�7����������g6�	P�g�:D]�jF��Hy�t�������������u��G�o��p���aR��]���7u#:r��5|���:�bp�ŬE�z������mu��0F�)G\|M�e51�g��m����3���o[�3/�랻���ͷg�^�s=>��=�O����������/���z��>|`!��r����;T� I��w��t)��#&��Or!;H��Lg���dt�٬��q8B�D�`Vя�2IKj#:�C0&�lW�"U�T�N��O[�BMZ��ݭ`g�+}7n�t_�z��{�Sy��]�Ƥ�Ν���7���_[�8R��US�����V�!�j�`"���o��᫾�k
�����L�	��7�����8Ĝ����gŽ�/���d��w;a����dZR��x��eSc����kX>������=��c,��e-�L< �����SK�/�˶O��?~��#7���>�߹}��F:�� �@����0w�7�n�����寞���ԕ�g����9�ըU��K�d��[���b<�q7��}�6E�q�+B�Q]�i��t�ē��(�܉�Ӌ�P%�:��]Ҏ��n��<Iu���OD������|�v[�k�s��w4.��g�X�q_6������B4㊇Y<;Ռ�ˑ#7�����,�J�.���շHkV�ƭ����+����о�M�p��O޹��ңw`R'��r��ā���3^��hc�ӧ��?���x���?�1��dm���ý�ؿ�����{M�bn��N��~ڥ3g��?w!���# �6KZ"*�
�ƶ���9�T�B��;K���A>� �"C@�w^��S���b�j��Dhy�fR��H��oٮ�7$GD���,��Q��vT&:��$�W��e�{ߜu��$Tҧ�t/2J�q��+��j�H���F�ǳ�ál�Y�@}T�������c�>�|1qMjh�)w%�U�:13���w�޳z��X�g#S6��L�*�[�7��� �w��מ��~�OT�Ld��"����h��d3�&��˱)b�Q��r|]R畩;����/�����S���O�m�|��<<�������0|��ӟ~iz���o�\������?�cͨ@G$yf-�q�K�Z��C�|�h�?�ư���/)�FD��|$�W����V��C��nx�w�S*�0��`�%_�(ґ�&W��]�ӧ��x ��ߪ�ģ���W~�`��>��������8����2��˦��F-�����|���k��kU���\0�9��J"+�[�n'�QSTM����u��W�2��O����4�������)=]�[�}��* 
p�^ރwf��OV��fvh�!�ď}qgys�O�f���>r��ҍ|8HO��c&�����|��.�^�ҍ��ϟ�\�5{I�ؿc+��h� ��JAߐY�a6��pQ��Z��$�3d��^$��3�l$'d��J��T�+m{���f:3�i��]HL�Uy����^>�'RK�����NĢ=��|6�l�c+G��XC~$֍/��/�e���%/��bd̪�$���U񅬆��c
| 5����V�=)WL�Fz��ɜ�v2:h, {&�1f�\Iaeß���uBS��ta�\��q�L��oA�ɿޥ�9ݪ��$���v�2Ѻ늩{��U����҇u��/-uI��u��v!+��8p��FއƛQ�&Z��X�,������}��Ɇ��0�ߖ���r��G�6�"�E>���W<e���?�Z9��O�8�"ڎ�{
Ѻsā���QK� ���B :e�뾈�u���� <��ż�!����K����K��Y@���C�I�Kc���7��~����S�F�	$=��bz'���!P�Yx@/�c�����L�R�^����^�����ۅ����۠W���V�^�՞�U�JH���R�s�+ߙ��{x��-��<]��&$���|U��$Iǳ�z�Y�2F*���#�mrh~~vcb~�������ڔ�UE~������b~ߞ��W~����^[�x㩓��`�XWX�T	����V���vk*��׆ i��k��0o���֦�+$�N�����e�\za!oļ�������W�z�^�`
֒^7k%�C�>��R!��7d�8Y_X4�k�8����eԱSgN� �0�`
S�/=7�I��߈��p滼{��꩗LГ���;�*�w~p-��4*��+8���iq����^~%�o�kKs�z^&�X�b�Z?t뭟~�����>z�����w�N�ϋ��|��֗ޱt`�;Ο~��# r �Iӆ0�O5
y�!�*�\�#H,�.�p���+�t�.�K��8�}��l.�Yߣ�\!T�����o�3�]��|]����l��ggx�6�w!���<Lа�aYN�n)��m̷���K7M:�.�TnjU��G�H<�G���ޘ�6^ة��V�����D��+������*�phR�������N���Rz�v[���S�J�P���/�6?{h�����QM�|̘��g<�kN����;!�� j@7�QsU,̑z�@��~D�o��W$J���Wi�����Y���&/i��iDH^tu����C^D�W��ؤ�P��nԈ�&eC���1Q�9�}+u�٪�F�b��=��R�t�+9�4J��w��#7d�Υ��rąem�\T���.:�1&{cd�jvz�'0Ի��`���װG�
�����z�c�!���T&5�Z�v����aΡ���A��[��QgzV��qYp�!/�S�
F9$��_$/g�onj�ݙ�[��6~>ƈQ��œ��1��g�����y蹵}A��Pk���P�{�p��|�
���uDt��Q���
����M�;�i Z�(    IDAT�A���z��Ȇ�$����J|���r��<��~�JJ���w��T����ʵ"G�����5n�6ÉI�:�ݷ���:^֕G�Q�]�����R���|�����/�o���U�����p��{5sv:��a��Io�y���v�1�hf\�^��鹩����55�I�'�$�>&�}��Ϻs��cߟ���ni�R�9��u��{e�G��8.i�M��ّ[�tŝq��i���l+MbW���k��"�����Q��J�Ew���mq\%F4qH��0��6�D|R��b�����+8��//s������e1_``*4Ѕ��8T��Wӝ��$t<�����_%���dV�[ƣk���ge�O�j\���GȢ�<-��~י|���~2UT���V�-d���&p�A\i�+[����ixe?5�rg{cnwfϹac���6e��D�����G�.^~S/�q~�;��f%{�	T�.	 ����p��&qB@i;"E���tfw�w?�;�����g/��?]�5¶�:L�)�Y+�����K��tkR��NiH�Z�������pI���]:eˣױ�������4B7��o���o���=2K��ǵa/��_�>�wX�������Ckߥ'0�(��峇8A�<�t-�>_��>z���{����?�l��E7�U7�RKn�F� �WƳ�{'N}+a�/[%1is�W������S�x^9N<�z���x�ίK�e�.ť�^7N�ҜU��!�t/I��Ҁ�RU�Ґ���t�M3��}��W�u��O���)#ϥς�b��!ӣ|{�������M`(sq��.��ΕOz��oD7������������|T�2UL�|`wSz�C��D��HeB�D����j�=��"�dƲ��#�%W�������/6V_nj]�p�h<K�5D^y'����<��Gs߉wm^��o����w��w�(N'��n����0��4=�o���u���¤������?~�������p~�`l�Wur�)ӕO����^�t��`�^���^�w�o��;�V'sgcF�{��\Z�A]����=C93;w����ot���uC�EܦZt�_AT��`�IZ-4X�v="��b녺e�~ @>���y׃wtY��`!]�|U�k'-�밺�!��i����Ο^��ʾx`xA��_@�_+�ʧ��I�OX����
BX������y9�<��奣��������o~�!q�K���в;����g�l)+���`+��J�ȧD�6s���~ol!n�t���Jp���粠U�������&�o@���7�ẙ;@lB�[ٚ`:�P ���u�"W(/n�<C|W�C>���G._z:��8�*XZYWผ�In��iy��c�������~�
~k
�Tp���T���_O���
�t؞(�eX�m��v��zW̗:=02�:�ۜ������I��No�@>�D+�.Nm�f��I���J}�1^�N\�����a}{����ŻS�Gt�^��j�[��|Tq�_˲�n8��xTP�F����Ō�B]�.V
�#f��t���g�]�B����ECZ�m���&I+�|��fr/���t�K�$��;���D�~$E�)kE���X�Ȋ��F ��2���K�$��a����^a�n�zW)1�7����a*o���O�ޣeyU�'��U�x����l�ٟ���m��2�e[�c'ZG~�3��~�r�ک�d�R[a0���][w
[�5llm!-�OV�e�#u�"�ɐ�s�{�O�$�u��qM�^��	]���Y����[m���3�8rլ#\����R��!@Iki�$�������/smp4�,Ď��oq��v�{�2�n���'ʣ�8�(#�5䤪t�6�+y���z��(���0����c#f�7y����i�{a�\��Bُd����'}�'�5�B$�ox���t�-�Ui�~{(��])[�w
���#���Rv���+��
�v����K��ܸ�a8������2���yt��<�,�+�?ȮB\1�HH�BР�������X�;QZ-���1+n>U�ѻ˙]s#N+3�b��E�� ��	-�����S����*n"y�ǳ��ӞG�I:娑 ������>W\>���c�	���*��Cj7f��
��Ԅ���ٟ7<�YώE&[��-��ٟ�%�4�C��U����?��/�Ҕ35|K\~9����邋N-�_�|HyW��\b���'S�痟��/�;��=����u���{� �<Q��^AxG���W$w#gϧ"��H�C/�?c"i�u���L�zz�����ǻg�����Ov��Fx�l*��\O�g��`e�k�ӌ��^�h��HZ�z�)�;��ӑI�<�7&=�0����o�NX_U4r8,;���re|����Oy�𲗼�xA>�eU!��tT_&o��{�bh�ǭ����w�v��<=w�0\"���$x���ލ������ B���s�v��Y��X�߉Ț&�tˍ�*���@�˱�D-;������t����F����� �'`R3��-Sl-JqE�*�Z�^�	2'R�PD�UR�Ce�Q�'{w1F�[�3�[g"׺/"��K�[A�).���u�[?�{�<�7��I�G��+��`+�_;�/��78��-~�"e[)c�n�")W�B��tɊ(�O>�;}����9ab-�3o�M����l5��j�疲�KV-e3���f�c�����d��ȅ=sSi�ᡝll������le]ힽ{v7&��H�'���q�φ [(�iE�0g&�;1��A����K6Y>ݭ��� ���p[��(����G��2���B���9'q�tյ��*�����yYjP)^��W���z�Ԧ���=���ɫ�W�8N�(]�Mcz����p���匿c�06�%��Y>�/��R��v����<o�b5��:���UY>��ʋ鱗+�1�U�����O(�I0+Z�VC`���?���w�}�����~�44�Hh��� 9N���K�-Z`�Q���C��U�{��W�5^N/�U=�8��"��s���|#���Kc���c7.�\�ɵ���/M����h�ַ�0���n�_�ɷ4��HW�IFI�]kWhЭR�5(X9`Q	U_i����#yE�,���(�3�����7����YN�83<���*Y�iVa7e�����q��;�=}�r/n�ά��	:�$�9����VM秪�F'T�2��y��?�j�ܽs��/�Zd�W�(� DjAL��;"X�ᣡ8�	�[�b��#0I�Gtj�@��������h%y	wm��������-��w��{��(mO��G�}�KO��Elq�o��iz���޳{ﮪ�(^�#RB��2{��3ّĘ�ۦ1�{3ҙ
��=V^����7�B����+��A�͑���޷��C����A�dJ��S�;���z����<t�(��v�&����uI�ai����LC�4��q�w��_u��qF FB�[ġs6_UJ|�5$f���(u]��nZWN	��o�����<�7I��z~y7�OF�p�W\���@Z6�|�1].�*1�/߄V7���Q.�6�V�eN�kJ��N__|m�h�ԓl��M�,���T�����zD*�z��g���������uE+��.���C4 [6鞼�?���[�!��2f�xs�������`0桊�-���8F��Ȏ�Y�=�?\}�	����
Na����r�� �E��Pg��w��7D��->?�&���ɧ�����z�^;�H�N��siE�_;�^uj�V��}1��}�?�P��5p����\�~8�zZq�{?y�|����ԇ����gy�����?���W�Doy4�vOj�te���ј�ѫ�Ԫ�ұ�����]��d9{S�{����I|���|�<.� ��[٣7E��Å���_���t��U��b^LӃ�l���k#��smU���z�'U��J�w��ܒ_&�Uy����d�sT���֍w$���t�t��x��2���7��Ǔ֯O�hT�e����W��wqFگ"]�/8���Xޏ�<��n}�Ϋ�/t����H$��$梃S;��7�r�����=ç��u��z��p�Y+�y�_���Ut���7?R;���B?�<����x��Zp��=�,i��!a"[q�15�5mj":C�$ ?a�Ȭ��I�^�2lڢ�v�t3]$� �*䏈�s��ǉ�5Jk�pa�+�������?ګ�������0~�߹��������޵?K/�x�=���ӈK��W^��}�Ucz�^�g��w�{�����y���w��S[���{�N�<�#��;L�����d��w�o+5&��7�0��>�t���I�Vf/ϵ���a�����'�V��������LF��%��޾�{��+i=Lv���H���uN+s(@�y��ԯ���AcBH�Ii������xR1��+�Qِ��	ʰ� N@�N�'Mu��ֶ;"/K�Ә�f�6���Z���	����R�*[�|���;q��
�U(�Ӌ+�n�F5������|*⺧�A �ŗǇx��b�.��=XG�;�f�>�t����/�����o��on�	;�]#�-��l��W>�S��G��*{��h�����@V'͆�eUJ��V^���~���[��o�R��~fI�5�-r����u1�����`۾�� �s��*P���>�|V�v�g��p��ϛrE(��z���ؒK��8�����`k3�b�c����d���Gq�OB�LCh�{:�́���K��^���myW�����\]>Bj���z��Cބ���j��J?V����B�{�O�1���W:��!.�VY�)sq�ۛ�����~�R�߯z��>�/����}�p�����~�6���~ș8Q˶��%�jS3�'��Өغ�2<���,ip�Sӳ�Lޝ�3���Ԥ�n����m�H2"r.�B��m+8r�8�I���"�c����b�D�-�c �{���þKmr!��!H�=G��<�G'�&����-�M>�#��廸���I�&)�=y������ڽ�͓�����j�����_�Yp��P�	L Ʋ����Vޣ��>�t�}�~��|\͕�ا�έ�ɉ8�|�K_:|Ƨ~��-����=<��o�v��_���ĩ�ɣ�䟊��9`�p8=��,0]�eñ���{���OfӚ��L�'
���'�>���3�eH��T�%t�}/���uƤN ���J*cdӿ����B���!��$4�F-�1��oN�9yY�W��?O�D�
�+X{�L�b&�UNoT�`y����������)�P�?J�����.�����O��Qo&8�@�D#_���UP}m:<}H�K��;ʂWe��.������k������A��S�����=ï��~��>�6�ptq�[�e'��ճӣ�������&��ԫ�0 K�o����(���h�_��.�^^>2�8s�� ���( �����}��	ө�|�y�
\Y^�s?��>�ޓb9@(V���oz��7�u��}�~���=o�ɟ��:�#,.�+��ʸ6�r��v�Gjh�z՗�hl����;�����lͭ����֒��	��E䗷)��1��Y_Á)��P��z�����^��ڜ�.��?tl����:#k|o~���[��IɰC�i�(<ZA���v&z�s����$2&FGA#��3��չ����z��/��jHg�س1���_�_;�c7
�������{���a*k)S䰖<���`l��q�F%�]㣚���S6b���'h��N��ر#�w?�  H�!oT��Ґ��g�7�rg݀mo����l~%vR�:G�����[*	؀�U�9s�B��;|�w|{�Nk���?�#����	���ј���{�a��ī�+��+r<�E`�����J��^�A>���J���l�:��-��]��L��ٟ��÷��簊?�?0��/����_���b����3_��_>�������2%��0�������3)-����*}7pe�y�q(=���՜t�/����������-�Z"~���_��_���0Ҝ*��8T�ip5H��aS�{ev!���q!0������1���ܟ(\��a�;)�rP8`��X@b{�:�L-���Ib._��_��E��d$�{2�0x���}��8>�s��q�)i��HC�k%�r�,�G��޵o޷oms����^���d�_�_P�Ol�Ԇ�V�W�o�=��՗���>)�`r�]���O��=�)���\��;���%a�����;���m��.���ۯ��a����ׇ���/̱#�~�~��%Y��K��8T�B}�O�upO
��Fk�|3=�י��gsϥXC��l���a��g�<8�����m��c1���b5Qi�/���S�����-��nY�S驯�b_�3�ʋ�ȝܰ���G>�3�m.޼���� Pq'�K+@���y>[��ǜǬ�mo{[I�8����˾,��;r��㱶L�|�wf�ǿ�3dXItϘ���.�3�z]A`�
9�k���B���g��q��|���~�T$;��E9�:�����g���\}���r�9�I�w��g�D�x��v��������C�E �x�;�#Y��ַ�%R}e������P��?"�_���}o�+Fcʿ�Q����v~A��u_-�����w���Y�n�������E�F��,g�:9�J�O<�p��7���Anػ�+���iП}cL �&��}�}oM�ϼz���7g	[�2"����?�����?�;<���°�BL����W�{@�Kna�U�+�>����4����>�6��ew�ts�4�o��?���I�?���5$�+~���3�п����YHW#�82�V�Y��&Tp ����XjFk�d=�Cf:i���Dv��xu�ո�y���Y7�gk�����#Q��ﾲ˷�H��h���3U�m��#=���O�VNb6��ȍ�2	b"d5�|=�g� ��I\sX�c9~��>0��������^�ۤ��^�d\�V�)����k���M{΁����Hە���4��Q/Wt��������<�T�O��ό��[�\j�C�X;������7���R��TK�Z���.��M�W�I #^�f!��ɩf`m� �r�>M-�IO,%�'�yjT���_��+�W����K0��6Z��A%��ظ��a�GI�d\H��*��_(�6�7���&6���w����_ĕ��ѸH��Bڨ����׿\5��J��,?ݾ2�{�Ǫ�>}�'>88�@5p�^V�zW������o=����ܻ
tp���A^��J6ݜK����|G�Ͼ��/��M�U��n��v��ʍ��F�ꃦ�VWe;5�۾�j=�|������f)o:rc�{Q���~���9��Ï�~�A�B��W���~���6r��Ɋ�$�.�I"=�������3��;�DǛ/(2:@4���>$Q2�,W��BN��� 9J<ibU�D>���v"Q>4<�O�@�͒=/Ӿ�rP�#a4�=�z�S���aLi���eԔ.�FnJ\�����[܂��`^�o�G���nd��/����_4���Q�W^Ș1��).�	�|V�c�gd+|@@���o��OPʋn]jNf�o�*������/���w��� ���k}��~�Wf&pf��_~Mj��z�R���
�wW�m�{Ե������
���c�Y>�s>o�_��Ұ��ON��3ܐ&��<���{�뻇;��$q^����4|��}M�ٟ���͎\�p���1� W�Oj�?��)\�sOM�9���r:�v��ԃ�x �k�u1���R�[�,q�}(=7 u��W��v�l�a��� KE&#-x���^R2���l�^��/zQ��㮝��Ï>�ٯ����1��e/)"p��������%��}5�Q��'C��i���=WL��c�����%1������J{��r��w���QJ�!����=�V��_��Q���    IDAT��n����+τE������ַ�e��O���<��#�Z�VQV?��O{Z��Ǉ��h���=�%��ww�R�w�F��O�Hh����j��v&����e�K�6��~��_��_�l��^=V�;I���oƔ/]�bXLj���P4��zFǏ4&ox$l���o�Lͦ��i��̮K-�0��r72?��|��g�����)M��*�Uӯ���Ga9�2{���
�Dc#G��w�n�P�|K0�I�\�<z�C�4"HZX̠o���n�0��$��BL�4%+����_ؽ~y�K���I&?g]�G�!y#�������� ,@ӿ�Ù�n�����Տ�*����dS�R�)��kȮ�<x
]��wy@X����g�}�;��[�7�H�����|ӑ�[n����� ��F�������B���58e���3�4h�0Q`h�a%0�&ϟ�@���kH��	�ӳ����������wxg�"t���i9é�xb.6�c����o	i�S㔎O`�(���[�ի,_��y���z8��1������ǎ�i��/.�wI���%v	٪� �Zu���c\���m���5*�;f�����
�Or�߈�@Lg��wI1�wo�C�u�a�~_0���gc�f]�?���CA��p!'<��廢,?>�$���<Z�1�ܫ�?���V��	�������W?�_�x���w�u4=ȥa#B���MpX�63�6i~����п�|!��j�,K��6�z�k��_�Aazk�&�^�������� �ıJ/F׆K�DW�xG��l�܋#(��zF��3�$5pV��|{��\s��ݙ�����(�!�I%�
��ݥ��{3=�ƞIdȃ�MDZ����$����gϓ`��ݩ0�ެ��Z�r�ﻟ��&r �#���LcVVkdm��۠���t�X!�8��m����{-�*ǩ��6b����[���x�x�.~T�b:����H�{ۼ=ߚ�.i6�A43�:a���������O��텃��c�|��7Ǔ���G�j��kJ�+�yO5�o�U���i��L�����>b��9ٍg�k^�K�'dy�������H5(0��� [����(匟sΧa4o��l����IŏB�Uc��O0eNN��(X��ӱ�go�ƶ5���듄���|�ȯ��dN#LcQ`�ӽ�]G�g��C�F���I �2C!�OB�=�:9$� ݴ�]��U{�a�K��A5/�2��_���3�,^�^Z$�j1e��^8�'V��4����P0X����\��-�{���v�v�mW'Gj8���=�B��oP�"(�4�*�Ӆ�Ue��Ry+��wo4�3k��yz^m1Yv�������a��/��r��+�\]<w��P����ϖ�O>�\'�6�ԊW8����N���A819��ẘ���ޭ�L~��v$�AGH� ��R�0F�f�1k��vk�Al���a�و`�ࣙ0�v�M��t����2X���ЧcT^#r�F��b�eOhAtG-���J3B2����Ԣ��at'�Y�D�Y>;�n�r���j6���9R�zT��p1ug;/�>_�m�U���I���xR��Y'�k�Pꍾ�#��<�0k<�K7��TX�@���icN��վ�[Z��<&g�ங �0<p5�쵿�_+�_~�_�A��	g�c������έ<=�\��g�Q*'|�� ~��Ō�0 �M��Z���a��y����#�6��O�����D�k�P�0ĐĐ��v�&���d�1�JBZ뮚����#�H)��FD�+���a�^�RMO�>dq�ԨEy����Y뗆���̬�����c�vG]��O�!Y��zzj��"����A��N��/�y�H�yO��t*�qL(a�����x���𑴘�`� ��#�yYL�Ӡ�.x�Ȯ�c���0��?u2L�E������ޙ�	������	�ݎ/Я��o��M���]Ϥ�r��0�Rz@y1���2�3����'�����mI��4PyD�f�Y��[�0Uë�\/s�����V��R �}T�=qi���:~�x!q&-�ַ�đL�$�_J�O��v�g�T��q�Xf�G�ϓ��j0�/	����g�K��0�l'`���{C�W�1�&�WVNֽ�9�Ue*�85&�4ճ$�Z�Rm�qb�|���V�_Q	��`���J����d���f7L ~����}����`�)��1��W�8a�8aϬn�\��ܘټA5�0#��;����lcv�C�P�E]�7e}$�F����z�a �F��H5>��b�:w�lᔰ��	�C�r͘�"��N���p���Kq�:Xyj �"�`�Z0��PL¢g����e�F$�n.̡�ui� h��fU���~v�������r����R'}h���r���v+]�pVSS�1WL99�f����AV@��L�t ���c<�Y\j��z��c��`�����5k
�|k8�BzoԞ��BL�9�0;��j��Y��1&k�ڪ���Az��O;))��.D�.=8���2��`����$(ݐ	��;��&{ab�$�3��BL��w����1IO�b\j���ķd'�����N�lG�۹��!�.�A��Ԑ�2�_T8�j1@��աzb[Dx9
�}SW?,����2w�ڞb�Sz��J���tS<ƴ��k����R�t�1Q6�2��z�jĭ�fT�d[��Șj�b��"Q.��Y�:������� ���ވY�Y���F1��ҿ��b���gWwe#6SJ�cV��-d�ާ3y����%�4��[i�lX�өMD�xQ�lS�<gZ����)��E@I��*����	�>�`Mo��*wz衪�S����g>�`�������^����/|�pv�����ǆ����j��;�R���A������.��}�{����>��k��b綀��WN�>QL�LkSL����=�����}[	*s'N>V����%�1<P�r��0��l7�l��o�3�.ޓ��e&�U�H����B���>�qS&N�<=����(�����a)���n
��I)]lx%z��X�F��'Y�]]=Y�l��t���H��O���*��Zx,���3��G�v��
o������i1�q!2���EV��S�ɳo�!ܖ6 �VF�.����$kҊs�B���F���	*�S��S��J���|�5�:�8����>��컟�n�3Ir!|S��^�Χ�5�-.7%_�tV"�����|�wg����yN�>�y睵��ƛ�S#�Ǘ��*�iO{F���;�|h8P�W8o��o��z�~�^l��mӱ5&�:V���?����w?�h��OzY���0�t䆚�����\p�n8�	y����^�&��Kʅ��~)0���C~��ǆ��W�Z�3?��´��i�ǆ;�s8u�԰�/� 1�Y��-�^mƒnM2c`L�`����U1��g�v����dH�9I��$��K_2�쥟8�IV������m�҅��h�!`N����gO�4�7�J����|�/��Sgn��yW'��`
���c2�M�O9]*H/���2����.u��}D����Y\��AI
?���q#L���X]��5asۭwd��=��T���bq���RU�?�̙S��q;��p+�"�9w���$�:i���f2O��PT+xbb����n���9|�wwԧ#Uz7zV�O�M@���I��#s��2�����
ZB b#�"����b�����~��|8��L�F�=�����с�y�~�
?���E|:"�4���0�3�۲�s�*�y�`{�b�0	��g�df<KQi0���^[?Q:���_;<��G�,M��A�����
�r�b>3��L'�_L�B �:73_y{��j��ܳ`·���Uo��M��̴"��7�T������9�	s^H=��L�K�������?y���[���Yׯ!�z뭥_����5�u�u�Z5e�e�|��B��p�L5���� q�\[�0�5�'3�R_*����U��\z�'N��i�c�@���p��7�a��8Y���M�&&2�N~��O�˗	����Gؔ�z�{j���}u�C
&!I� I�id�� h3�����vt��<���ܘD���F��d�0dC`�+�8yr;�a��(}/�l��
.Fb�o�Yg����K�=�k`��w?>�|��B�z����s�f(��ԏT�ٳg�T
s�O���~�=��c�d0����Ԭ���յ0��Rl�Yf�05�y��ß��ñ>Tyr�GT���OD�&�KÝ�5[H�������^u�!%�L"Tc��v2,��m���a��c�c,�y�*377�0<����>������|K��&��L�W�w��a��2��c��58 3:����ܡ���L$��f,2Q7W�Ŭ���O��O6S�0��Ӳ˙�<�S��f����_��V��=q�^�����B����Ioq�'b��$��*L��Ku�Z�g�DT�)]1�kS=�L/�"�B�1&U�1'!쾬�DdV L�����՘�$x�Ɋ ����������X����E�5d��a
�D�+K�	����S78 �r���b�L��iې��Vd��'C^������r[�Nx��fq���A���ΕݚiV.?��psq9k #,8�	ǎ+�'�-q3)$?*��oU��.u�3p����'�����	�(��⻸,7`�&���F���1�vUN����S[f��?���/^<�>�53a�0r�~Uwڐ���|w}i��=t��0����������
!,�N<^����ʦ?�]=z$��ܼu�����~w��x]嫬�GW���S�����t�✄�{�J�3M�%	�2��0K����h��9q�������VT��M��3l�$]��f:��8�pC,� �<u���O�����	ʜ���!]cYy�Ր�"=S�����P�'X1�c�Ϥ�2HSf�}�3xNc=x�p5v3��F�iu����6���s�:��n�%>�Hp���Y��[�{�bNHH#W>:����Jo���*��2���䙛�W?+�>R�.涅���r�^�VP�� P8)֥���NLGVo?��O����Z�S�.� K7'YI)W�R&��1"�=�<�NBC�r��Cplj�lka�!T9�0�U<��}������M�THM�N8�����1��+���"�y~^�Z�"�M`�><���C�c�b۾AY�Y�M�M�I�;����&❧̩H��b-��9H�KM+c0�:�^������}	��|�����{��b4�o���LV5S���͜QC��Ou1w�̰�ṉ覎v4���{���C<���������=�2��~�a�������]����b�7Gv_<���@���j xf��G��Y�2vlf�w����^�BI�t���|����0�9�WQ�^��7{��/�[/�N�,8	]��g�6������E7�0G^���������V�X���%SFc�ѻ�DP��`^�k�>4.�����Rl��PK�OT_\��zZ	&����~G� ~���a�e�&��'��_��:j `0}�`R8kj�P=���^���翨����_��eW*+_���>�V>��\,A�(���E���ތ!�1/F孨�幩���6�s=v�ԯ��l��<kϓ4ДcH��Z�����\ a��U�<�q����O�8\s=zr��Cޯ�|d���X��u~f�>���0]�u���t*����}1E�I:�F��W��R轅|1%D����`�����.+�4�7��ߟ��%/yI�ʚ�f��^�3y������/���_�6�� 9ԃٽI�b�b����YPV�O�=O:0��l����Ņ���ȏ=�h��ʛ���{���(�U0��$�;���b��0����\$��}����V>�Y��A<�`�)1k*�L�p���5B��exzWw����m=�ͷ�:|𡇇W}ŗ-^��7V>�}񈑣�\�9�����<]s�&_,^ԁ��*e&Np)BE�DBc:8S�*ݺ�6���xf�N�j�'�"�H��$�쳚:̼�U���n!p1�w�nÌh�]#{�A�Z#�I|���_��@��w����z�ɟ�ɕO�@@�ӹ��2��ꩧ�^Μ8Y�l��d�88���f�FIKRo������E�^��G]����G�_
�F��t�r�fq���Ï{�[|²4:7fꖝ?���n����?���q%�)x�F{o$�Ñ�}�,�/Ʈk���tڢ�F�h\wá���_�=�|;��o&q�LzDuRi5���AF|{|ː*�t�1�4�F�c��b�cY�s��O����bHa.@���d��Fæ�U�W��K�U\����ڥ b4LAo�������ݧt�G�g���f��L�]�|L���e�|����<z\���`\�O~�X��&��V����Itp=�YϪ<xIH�/3Qp	w���;+ǽ�� ��]/�������T<��m���o��o��"8�f�/�@�s���7ɣ�r���{۱y/�G|���׷����;
�˼����H��pUpnց�����.%��RI�{��jW��������piĺū�@*���\'$�"q!B0;FAqUA߼��P� ��!A����xؚ/��aqC��cV�>�"6�)��\��������m��1I�$�;1KF^E5��I�ybd0��� a
���l 	�Sy��lM��D��q��b�^����|����/oD�_ǗzHיJcg�aF�wy��3���wS3��~���C��O�W�C����|�(̽g���+����NX��Q�$`#@�O�~��pU�<���:ea'�M�iѓO���p]�[�ssM�Z����R � ��š{A�{��'���Ge�w���U� 2奭HG�b�*?i<K��}^�꾥GX����퓢�NT��y'/��8|򐯺�/o�XC�W7���=�I�����m8j�>l^��Ă!O����,Nz�p ����\BY\�+��dA�^�Ա�ȇ����~�d���p�'��W/:�{0�]\�$���w�������#�F6��$��D<K����ٕl*㣒��~�n枞ܳBʙ�:x�@DBE��0�4��j��qk��@*���a'�	f�*KM�T�X\�e|�ffS>��Uq��)��y�-e�����
LZ`w/�l����IR��R�}�O�W6b�N��ʛXjvh������V6��[�:&��K>�3���w��3\��[�n�!���Jg6�@�����\z(*ޅKm���R	�0+�EP�^�p��}���7�T�h
�u�my�$wT2��+�oG�c����l�ds����Ԗ-��L�GՉ ��}7����B�]v㬅�?L%ﺙ;��A�M*kUղ�PHѢ1t�g>�9�'}�'U7D�k�dIX��b&?�c@f�)��o��o�Al��=��YX
8"�f���ַ2�M5k��;ߥ���㝠���it1V�&�|G������`$!)���Oy�]]2X�Ay���3��g�E˳M^�W���Yj �I孭���`J\��:q��W[l*�:;�L��H�����{S�ʿU��-l�4�u'ܔ)�{��N�i������|Wwxڌ��_TO���V>���]Y�X�Ѷ	���?���6�XP���~���mA-&aM�k��(��1{]�T�p�D��>*ܙC~;;�X-�t��Dب�،-z@8:,�ihn���1�]̔9	a1�[H���������Ǉ����wv�W��6-i�ک)�V�Dz!�ɓ���
�w/�Ęm9����F����KM�PW�~0%��zw.�򭺏��덾w�]́CL���1R����@wT���27��_�,��C��y���9e��Jởr��d~��ձ�%�y���3ñ��m�V0ƹ�Y�p�    IDATtq�E�[Io2��g"������DE����Z;u~�;D��C�tԃ��B_  A�tT�k�g|�gTe�O� l������&����@=���]�3�X����x��|�^��1-��@1���>M���ǤHغ`�p��>'�tZu��ީS�)���
�3��OY��{
i���k�]����MYʁg��h�SO���x�[���o��֞�C���ys�M��mo�����&��� .���{�a[Yd`������pZ��Qm=�7���X��wzo����%w��c��`�T̢p�X�Ŭ|���l;�=��k_��2O5�Dwm*�Jw�v�L��A�!D@Jy�ePF��C�b֡1'k ����-�p����7���n$g:�N� n����� b ��4&=�qkWV�	�p��y���ş�3�̅���Fm�6&�Z���@�Q�J�gp#��˦�� ~y�C��5ƄRW#�D]0��0K�C��&T����y��G8�=F���i"�L��S��z�%DF�tu�'8��5�&�¨�6N[�	q-��ؕ &���튛�U��&�o���%yL��[��$�Ǐ��-_�0U�	!��Co���AtSMvK�
	�G�����OG�4ߕԇiH̋ M�kcn��ʦ�RH�4�"*�aj�9?U'��4�λ�1R���a4V�w������\fW`x�N��d���*����3��{��Ge	��=�z�y�'��i��Q���]���=�Й<��"5�Ӱ|�HZ.z0x���3���k�N�h�<�盲HO�~����W�Hs���6�,��7X�0}`�Ѻ�wfӝ�����~��p#dv�\�6������^�Ե�eTN�rl�fT�������'Δ]���bOv�Bx1�R�H����2<�݉�*�Ņ�u�͍9�s9��>��>$5G��3a�������;O�ܔ��V�Ӹb	����|n1z�v$H�Do_�
3MD�υq�3���Ҫ��w�b�*ͬ9�}���po�b�����-/ݜ�"&e�հS�]l�N��l=B�Pl�f�Y0̠S���~�������`�Č؊:d��a2�;����0��fEL~���7���a��N�������`�.�g�ٔ�8��l��R����q�8��̩�l� ��x4n���HW{��/d�k�F������Mo��o$co��>4���?��GR����lK���L�"�H��R�)�H�npk���嬄��B�����[��i��Pҵէ�9>��8��"�쇇&^>��G�&��,�!i!���V�֟��Mri�Z&����Z�����F�)�߿�67S.��8̍�+�Q!��NV�H/_�%(�3���9�I���H(� +EF	׶\$O�ϑ,8eq�$��J�Eˋ�3�"7�v�ӳ�<;��t|];�-�8{��HJ6��V���y*`U��R��A*���3���
|�j����r���,�=w}cex�3��_V�\<W�� y+S��b�V�=:}t�>&��=�sa�H��������)K�Ƽ��v�ܩ�jȔ��JJ��e*����u.��_V@�id��h&W=��Ne@I��c���9����@ʣ�{��ѹ�{��H������f�z(��?H�?\/W�R9KU��S� �!�F���=�����ѧ���Q7���m���b���_�j�H%�Ę&u� f)��u��?�Aˁ}\U�{�Y�ɔ�N��EB��J��H-Ʀ�|�me�Y[��1GE���b�\٬|''V�^�g0�6Mn�Xوq!V��Y�Y*@V������]ԣZd�!n�����:�;��f���CK�5���~6W�~���b����9�6��x.���d��?�W�7�t} T7�=Aؼ���Yw&�s`x��4��e�赳�fz���Y����l|y���ИW��pg�w>4�K���2� wzo���=�3LM-��9�{���|�~=�v2��O��������CZ����a�ލ ��
���5���g4NZ�	<��q���.w������/�/rH��u��Ȉ�F�=Db|2�x�U�w��rq1��L��ed��^��Ft&D��K.�dƴI��ߎ��3�E�u���I��ﺷ�˂i
��)y$ݷ�51���
�z�ɤ�SҒi�nX����ұ��xs<�߅0��ӏş�Ψ"���I`��
���G������Q� v/0��RlõΞS�-&̪&��=qӊf'k��ѧ�����Q�Dz�Y"øi:��	�R�4�������۲��7.~YH��x������O�F!��=��͹���^?sOd,c"�*љ
��r6���~����mk��l}{`1�	�=xv2Q>:�=�����k2-�:���0� #(_Pfop���HI��@���4���a��mne����t��?�>s����ax�;ޞn�^})=J,9�g7���3y�wbVz�K��P����I�+G�ə0VtPD�@��&]0\5�FOc�ы��@=㖭����s�3֘�}���X�Ƕ����$��]	zШ�a\� �@Ofܠ+tf�X����gQ�,�)t��{"���3�bf��H���8r|������S��o"�e	�����L&C��/�˧��؊��L�;s�ԥv�M���wT_��9�+@()i� P�u�C�F] ��j����./>0�Kr4>�����~c|��L�o�?��h���6<r��4��OR�Z�Vq倥36��,
�6XL����</^��i�s��������E%��r�+�gx��o�r�����F;YW9��#�2��������i&:����$sr˗����0�D5x�4+�2pԣY�y˭7�w�T����ca�>g�!��,ڥ����o�:�K��q�ʇ�Vf�4F���Zޙ�G?��;�Q�0	�{�k�Yaz�jzF��O�e8�	����vr�S�>;���s��إ3�1�Mdq���[����h	�R%m���ۓί'�O�/�G�u>�#��ѹ�����~t8�K��f�T'���R�ŀK٤e%��\*�E��]�����GO�S�}0*E���d͆9����{�D������".y"b�ЧtK�tx�@��I
#�6�� ��/=��lu��t���><��E�=~��񙅽s+K7<����qx�����v��n�	j{`k�o���������6]c���$4;�r16ɮ�!�3V/�������v����h3�5�Lfm�Dc��>�y�3��{�}-�w�+�̰C�97U�0N��a[ωR��=��F��e�͑M�~�'~������Xh���SqZ�f�'��>t��`9��U֨g�	�24,o���ն�����R5yAR}�ę6��-}#�/�~��X��0\�Zd�>�c+N�Y�ވ�~$��	Y�#$�hV�<ЛuM�#=�h[Ic�IȽ+�Ҟ��g�$u�R������p����|��F�R7Ds���Ƞ��T����y&a���t�`y����3x�i�$Ji
m�Ù����Φ+����ٽ3{�9wr���S�-��4��7�r��I򪃺��#r1Ts��}ߌz��7����1��O8�RQi�nW����2���'>e�=)n+����'����ު{I���Pp/�ш0�F�7{���ѯ2��Vgz3�S!�3مц�`)�V���r���s��Cs1�M�ʼ�������G���<s�Ԥ��3��6����#ێ���d��YK�Ӷԁ>p7c�ë�N�����c�{����f�">�����̗��\->�U��!�$�.2��
Bd���䱱�NY����}�Y�[����k'O��̆/��A{h�-R3�ɟoFR6��K��*�_��e��7�DX�Wc��㫑�����Z]����H�Ŵq!��}ss�1�/�LxaJ̠q�I��^���������~�NoC�JRS�����=9*�9�l,�ؿϞ9�squ*�'�28���icnj���ō�?p�o}k&B�H8���p15�Lo�5&7���z"�z�7���F�+��YF��4�e��2p�{ە��?�����K۟��>�'N<~8{�L�p�fj���n�p���Bή�>���GP4̠9��Wd�2���O��g`xE�k��f�9gH�j�1� yl��mE�9���G�sf4"_�����k���Z��	 a��)h�����	�����%�r�Y��)*jCt�c��0�!�gG?/�-,��ܾ�ӳ7�tˑ�CSQO�]f<HBL���<I�����2#���ZE�q6���w��$�%P��e	J_��'Oon�.-�lLL�Lf����ٹ��{������x��K*v\����t�Hs�2i�z�Dj�SzyI�H'�6`�7ͼ)�9wv}n{ϙ�3�1�������'w�N�n�D�����֞L�M��H
k�;�'���C���춘C�G*�l7���>&���+��]��̧�΅�&�{�o,��ؙ�Iٿmfyssgn+�O�XTM��0&-���d�2:���@�����Yi�.i6ih`�j�>뛗67���OrOl���g��������z�0MB��*u�,��X0�k�tS*�XEUx2�h]8��mtm�<4����,q#߶S�����w��C�fl�v�"1�.E�f�)/���P��U.�8A
e��6��t��0���T~f�2�����p�m���^��mN�m�Y?������d�:рL�'�1S�HP'x���`���tpfѭt�'�4L���0?+�U"xY�Z߼0�x`}'{O�]�ܘ�[����{�칋w�F߿�HA��z���5��&s0�F�lF
ܙ����D��M=���5�g;��&h+Ri���Vv��$��wi�dTǙ����'�/\���[/��l��,]�w��W�^+p���|VU�����1��3���qqq��㦓S�B���$�'����8����!�y�����`y|C�J���&D�����6��:S�p���M�ܺ���?k�#7]���_��޳y��O;��Ox~I|]�AZ�!䍉����m��	�����nNC@t0�8q���F3"�b��{��ژ|���΃�k;��V'Xߞ|8��^HCٱ�K��h�=�<�ԙ�;��x,��ݲ�l�A=~_��QA6�m��>�|~����2�����(��֧c�����/�용��sv�
>���-Ѕ<���ԡ�Ϣ>.?���]:��V�������KS{�]�
+��{��ت�9(K|�k�)�\Fw�v�#�\�b`h�Z9�H��W�6�� ���������}��-��0�}�5�K���!� ���������`Ez��fPi^����)�߰6�pxmz����ҁ�#�=���LMo����̜��B"�� {|L�!)��HF��b�R>�$���\�'\^�=��6������k'�6���{b~~��lTp`F�s�i7���z����I���3��&�U����yHc��u�ңŤ~a��օ����m=�j<x!������޽ϲM[��V�0S�f�+�1X���%e4����ϺJ�Jo��?*�Y:LP�� ���,e��g�7^��l"�ށr#s��[ۓ���Μ���3�͚�� Rwu�wM��'p"�$*A���i&-�E�d���I=��'��\��/�NI `p��жPݲ����&4$v�7�}]%�?��U$��p�\Xv>�=��V���,�GzڰᔣA�À���ș�C4pv&��Q������յp���nz�͜��_�ޞ٘��<�g��b�&Y�fg�lӋ�����5fV6GT0�jp5PJ#�p�+���tM����9Vzeckw{*:mN$Y���z$��F�S�/�L�xF\f4S�2<c� ��Z(�,G|��l��	&[����z����<�F m��~��]nw6�?���/��5җ�VT#�*���p��P�{�\�C;0g�"O�k� �5�c��+�.�6��[�%�I;Ƃ�w�=�xf����uUwC�4q\uO2sy�wn��n����͘��Pj6JyVi�>��\V��:5�!F!:� ��w��t�9�C�Mg �j�L�ą�.]��{�衻�3K�w&��9usb{����|���}WO�>���ѣk$����:B���O�~�zf�^����2�8�0O]#ť�PrIqM�]�ڝ�>�y��I[�]�!�s;��/d�l�`^j�C9�u�QM��P���x�iO�k��o��{�ynImh��ɴ�)���{k	O����}γm|��ęǟ����s��#/\�p��˧�w��cύJ��^�o�:���4��^������z `�<��5��iqa�̥���q'��AO��Z�鹷����_����s�V^F�|���F��ٔU���~�g�$�V����񇫲��K�]��m����;9�";�nf�y��w�Ο={0�*�:}j>��5�������)�H��#S�����a��k����،����F��_�ar��-7�\�V��.̬onN���w{hyl����e�S�졝��ǚ2��w�k.<��&m����w�1r]�}�;w��{���7)R�$S�]S�,)N�q�T�0M�p[@MӨ�?-�4(� h�(��H[5i���Ӱv�(�r�Rd�R���II+r�%�=�;s���s�^�bH�"��V�^i8����������A��kQf�@|6�駟NLN�H���|����f�TX|Y��<s]ŚpŶ�:�-j���R�r��6�7��di���ā��X#z�R�R�<Qh&����hK	f��{����}��g�]�w�L�<��(+�1Y����Ɓl~�c�-{����6�0a�z�x���M�5k���$"�S��㮻�2 ���W�b�
p����#��J8lZ�	�?R��[��`M!{43x�?w��333�v*[�����Lk
JP�e�f$3.�� �۶�+�T}�≉Y&+*A�e�-*�yQ1?=s�Tz���>2L1u�������u�ًsBL�m�`mRb�ǶL�vY���2�9dâ�s�,�����%m�R��._�|��E�2�׼��{�'ƚ��.z��۽�C�VUe��m��s���FǶ����d��������Ǹ�ey�Ȫ�Jg�)��#O��_K��ֱl��N��.�:h�����.-�	{0~ Š�r�};�O�.�-"�^��蔇�ؘ�V{ep��6Zu�-	��	������tqr����?��W��+ SX�_�N�W�.'��8pŲ�d�.����ժ����x��iYX$Fh�iwmɲ�Rc _��2
��z��:l�h]Qq��H-5ț�\v�=?��x饗_���6�7�F���o��9�%���w��O��jd/�l�8}��#�ꝼ��٩;v�=}���f�C����"W�쌡ZP3dbX�7*Vν8���[��8�de�:yR ��w���I�ڔN�.��fd�IcWd~� ��S���g����QˊmB@�����|�TP�P��*�R�R��vT��qT|'_�9�e��G����<s��lO�K�U�v���Vl��^����?��ta�B�M��{`!��}(7A�
C���(�j�mݚ�0}:�Ƨ�)�Zd�K�ۍv�z=){��gX:mUJ���7ҟ�X��X/���Û��2���ވ�;�i�-�	����+`	D�g��R��'�k�&��ʘ��X_�M2��@Q�e���*�,��X�d��̅}A��r���7ҹ�����z�����}�*�����?���c�^�3&��xO��.,�*��v�#�`�>\D�  �l�Vm(�� ��P�h[����/��WYJ$��l��BJY�8�@ 2?��(�  @f����I���Hjm�<��c^��.y���pə�T/m��=��� "��X[Pt�X�i�)Bn�FQ
�����AQ�oY#�g>��9�W�YW����K�)9dp�P,�N6����;�n��Gg���Q��    IDAT�JF��ܸ"d��������|簢7˦�{�>�U�wH���Fkc��9�C��_d�����p{�7����E��r9������l�zǏ�,�?�䟵Bnco����{�wpq�U� �H��2?iU������w ,@ @E��+5a������}�8wN�r�8 @3��4����b��k��`L�� �g��Ŧ�)<�Hy��/�ӣ���G�w����.^��k�Zbt �k5Ŗ6��6D\�ܓ{�"K���8
�N�I�p@0� ��.s�C��4�N�h��rgK)i�L��Rٿ��=��xr�9�֥�Sw%J��c۶ٱ�b�8�I'�6Wl;۶;�����~é˺����c��f<����p�+Nx�
m�ѽ����(�6�Qz=��^\(DE�$�(�EB�;hL d}~��o:�x�_�X��������`��`3�O����6�H���f�k�3s�;�p)��i�{��#+��t��9Nw���YQ9H��v�J[� H��}3#J�󹴘�0to�$H^غuQ���6Z8d�����`�Lt��{*T��te�˱��	�}zuzЛh�N�y�<!��m&[���A���J�%�&��
�	a]��.M�#;LD�~^�]�=�y�jZ�lo��쩩����cJ���M�_%��x���ux��P������a��"�p��T=�(wϤ�n~=i�u�`u�`�NJ��/
��؁[�x��$�}�aa;yU��Rb��5����9Am�{]��Sf{]tI�b�� �{����ų�����$^_yC���f��UC���2�������:j��M�@Mp���̄�rɍ$9�IQ��xrp���tUP��G�PTU�VF�'��r��d(�!�p`�q�2bH�9CV�!x�.���Z$�AA1����L*�<(|Zb�>�)�X���:�F���җW�*�.��WBW� n�ƹ�7Kg�׆C��A�%X� �p7ZLL�Ʋ.�97jz6mjdit҆��u�����n~`~�P�������Р�g=O�p� }�3�ub��#��m�1�,x�M)��M��
�b���1y�
ղI�G7�L��.\�f3���SNJw�s#%��2o.��P���^��1P	�l�֩���Y�(�^w7�#�֕F$�_ή$N��{�R�.�T�J̠I;�x��y�եlſ9�5�j�������;����0�%B�zh��f����|�K�7M��jH6Y�Y"�XG�#ѹ?�ތy��D�
�e�k�����S�A4�J�)BeQf��z�!����������4�1X�کzB�g��\����-d��a	H�G�@�8u;������OHi<G���B�?V����6��D/GQ%|�	�*]N��P,j!�D��f��/r�1�鹚�;$�aa�nا��� ���t�C�����<@��a� ���ǔ�����D�xvv��K�b�����>��
�\-��4\��5������ {C�!�D�Q=B�W	�T:2QD��o����o�[O=�({+ǲ��k�~.�x�ƣ~����f��V2�`@��7�l��%������s(��z���n�.0�ٝ<�+��״�=`\��W�57?����%�e�l4S���~0"��ZX̜77F >��BOb.75���]��{���T��~UhVFq�d�R t֑�)�*3��c�U��0��uQdE���1��ڵ/�C� �IU#�gg*A#��K�� �-?V�L�&�5�"�2P�D��X˟6u��.s^�"5\[شS~���_���Rb���,H�fT,�`���!�x�O3Iw����Gr6�3$8|��D������`�!�N̏�(�������n6{2���J���!5S!NOh�Ta-��o����u�������
��[X��?۸�~啖 �k�[2i<P�̂V��<G��K��É5���FHǲ>&Q���u0�G�BE���X��Ua�f5��#|������}��Pa� �n�}�/�u|�2��[\t��O9&O&�+Lhd���rH��\���'�AX���n�k�5ĆB���g2M�[~� �a�qy��.c�����A g���������̉q��^?	�.oYBe#�O^0��_8�m7ܗ��ۦ���K53-^2�`��$1�M���M�w��\ψ����qect�䝤�i��}۳�@��r��ي��c/��C�/���o���n��5�\hТm8C��A&2i���tEi"���ʠ%���>��b��~6H�`@����.y�ة�d�n�<B{�攊9��Hb�@iS��C)�l���R���Ur����a�{B�ru�����K�H�0�*띃;<���۩���K�o�6َa�8�I�[����/����y����B���y;����QOM�t8�i��/I?k6�K�BXb�$Q�զ����tb�
]
�)���Z3>8�6�o�aV/�Ŋf���2kB�Æ�c��k|��մ,ސwR��$
���<�l���M^���cS��)�t�㎛g.�!D��o4�-m�%�!�d˃v0v�X�v},��1H��1!1uN{���>G�tz|Zp��<4�ۤ�t˞h�(�;�J��P�&>�F���1��m4�$l��2M�%�)��*J���\�&^˱��*Tk
"&Eޙ%L���u`z�;j�����	��SFQ��ˌ=XK�b��������2XM�a���$5!�jd!�Y��0	�jޓ���>�������J��W��;���7TD7����!���������P.��f���T�(ϷE}��t^�>C�����zG�pȭ���z��/�_4\s�R�hqD�,���A�ɞ�(���-뙨�����0�0&e�2���a�P��Ź*�dQJfy����_
z{�)�z) ���=V�+���U�Q(��Tsّ=\����ƂsLP� ��%�Bq't�Y���|�q���6��|���o2�.l ��ńQ��V���`��޳"3:�p�m�W�m��%_h�x�����xB�H}�ėT)`��r�2��wD��a�5z-��W����-��mG��YM5*���Gbd�zA�����JU]���C�c7����;ClXV��͎��6_�+�n��[�A��l涡$mh��6e�v�|*,��::��\��`+�|[��R����:d��Tn8�"�?B�#SddZA�^A*�( Xp��rQEv`���5�2 dBt��"�w�.:b�8(#�m/8�E�
M�H#G����I���*�b�� �(�^nͭ/-�(����yR	 ?�yҝ>��Q?�w����B�I187:�e�>���mE3 S Z��k K�2`��k��p�akBI��1�k����EVmO�\#gO�/��83��͇�a���m8I�y�̔�.���Ի�'�d����8��5̣�0S�ծ�������Ξ�Dz��v����ʽ�	Kus+�Aq�'',�Jbp\!e���i�W^J��(��ӦI�ע�F��4��9+��F
aO�jQ7��W!��:�yf�$i�S�πQ��2�Y��hk���U�QY��A�����6[y-����0Y�^ngK��<�G�+
+%N�a/�w�)O����fՂ�L��*����G��>%)>�V�ƆjFm�o@���˱��'�j�є�t8������A�z���]�-q�L*Ng$���@J���y�3-���l��pD�e������Q��CiӲ�C�9�W`'��l���y�-r�����2hEa ��|��6v|�S��tU�-���uܢ���v�U9��H�hP�7�4B��1t�(̈`��.�I>���ݶ5�x�2�w�ni�<��`T�vғE�TSi'�;�2��1r���uS�S\�.r4�R�~��+GA2����@����ܽ�2`�����v�R��'T6�β�[�:⻪�x��BN*@g��Q�|:���Cd$�w#l�zC��n�������Ae��D��(����$b����	�&5��*ϋ[-&CK�W^%Ï4�-�a�0�^��`���d (�MON�;�n��6���ޯk�Φ�U^C@��q��2s�2��7s�;'�#֒�܂���|��|đ����ոu���u�Xb��i�+}]e�=B�Ș7�H�)|���*���S��=�oz��~rdr��kkUo���TJ����T_�1�d��M5�Ũ��ͷ���$�`ձNg��xz��!p��U��,�Q�v^Fr=Re�%-��G�]Z��/kguX����=��'�����e��U��9y��u�)���	pQ�Z��L�0��tt=lo$�[�ʳ�;����`=l=���f�jX�aOHՇϓ"Bb�z���w�[R~3}'�NvL^QjMf��lD�Ɗ
��Ϣ��r�4�i��}�d�`�r��~a��U��)��V9�i�qy�5�R=R�+q�ɻ�ʹߠaW�)̙Ħ�{�W�H���	���\q�3�K��~n�E��-2����:[�H_1Dוt����������"�ܥC�ʪ�[���.H;��x͵���$�����;d3��u'�rhA�;+mwtO9Kj�F#_�b'�/�dN��X�m.JK�B�Ѧ�[�]]qM����]�1��̷���8*����oᯀ��7���lT%>	��1m���V�%��y�&������"m<>ː�Ȕ�!~�ȷ=�����+��
w�D�����KZ����6l@�F&%�4��N�J���T��b?��ߏ���Z�J;�wۢg�+�D�7�U�%BN�7hg"�и�իfXݲ�����x�EC+�}����sK��(S��N?���߽�p
+��%�x߰��ˇ>I���Ŭ�΋GE���{y�.�'�'����v��g;����R~-�9�Ju���@ֈG�&��] ��q�I�[���Pǡՙ%t��j�0�'n�W�cK}U�.�06�PwT�ڽky�5�O�+^��TMϖ�Ï^w�Nl@�ɾ^�j?����<Q����*�8Sã���~��d��c��;��M�������G5����r�p�ͬ}��~�~�Ԟ�z����3e�spF�Jmz����')בd�Zʒ�@��Ƌ�s�d:!�/��5�}��g����nvH������;�	�n
9����e��bڴ����#M6(a��K�F��{BJ"������T����bn0���a�[�M�仝���f\eemI��K��p� ��Q �³P-BKfL�B	Zÿ ٲ���8;�]2�m;W��n\K�RQY_�R"�p�Jy�w5��(���F�+WO|�5\r��1���l�E�Y2���^܇�`�F��ʠ2�:a�/��jR��m�T-�cV�(�@�Ռ�s�������f�C�_�"-�a���.������J�'�Q�MԴf�<hPS �W�P�ǧ���O��v�^}���J;.-�>��G�y���Y�H�{��#o��3�D��ɫة̫F�6)��$����*�vuT��j����5$f�5C33�&;󚙝�)R~HA!�'cf0I˨�J�ȔT�����v�o���x �@�YHa��f����.�O������k���<���L�,N��l��lI���j�>l��*���.���	�� ����0��Ի����C�6:��ki>�"��ע�[cCM0Aň�6�`�,��Mm��D�dx�K$M��&d�*E�w]K�K޹"yL��5n[ʌ��A6����+�� P���-�q�6h���4�I��ج5�'�=�&@o�U��y��DLB������;��:o7m�����o~�F�C�,�,�B
>ྌ����,�%al�e�����r��څ��?#考̯�=Ws����d����%�BO�_�OM��ë���K��6�����5兓�$�Y��_�c���;S2Ȱ4�7�s�/ȣ���IS���dx/d���v�H��R�H�F^���0V��ȏ�w`M����cF�`Y�C��\n>y����>j�,¼��8X4�QE�Cĥ8֛H;WZ	?I!@~x�8��F\�\M]u��`]T�o;P:�0��yE�d���|rĘ�� ��_��]40]\���.�ktO1,��, ����k/P1@�m��:�K�`
Ҁ��B��
M��b3|�v��,���΋���4�D!��F!|����6�pza\�%E���l�i�$U8D�Kϥ*���<d��Ҩ���nD-aRwE�.7aƏp�����{Z~8P_�ľ��N���B�b��品�B���a���L���ז�(�s-n�aK`��B���8j<E��Z���בJ	������	�%��﭂U�u�<�|?�bz�#��v�?>r����MA���[~;�K�
�m�p��3a�k�̬*6���l�oJW�n���=:;Ҵ�p�Hb�5�kw3?�U���ዳ�$��7�M�j'�q���vȚ��Ӧ�#Zz3>�L���$
��
�[��&7��E$��鐺ο�1����̠��b�����]\��'Us��/�ش3�DM���4�_m�M1��*� Qw~g����n{��ɪ�y���Ǚ��u�L�҄ȣ�G��Sn,5ÚX�s�_�r�dbmӗ:�x�6������'~+����Г���LU�.]�{Ԉ����h����j@����'�.y��x~�	_����MAsñ�6�<�o.�??+���Z� l����l/��R 
_�1.��x��ݤ��bVM,��Ҧ�} {�yi����+w-J:��'ko�|��#i,�j�8���qfhn��h�ٓ�Ԭ�{�a@B� �F�e
6Y Y��̷W�^��~�R3��St�M�Ɇ	z}�jw�aG[	_0+O����@0I��ק��Co-��X$ĵó�G�������?���d�"5�R�3�1�����ӑ�@��Y(��j�'4��	����@3(^bܕt��'qC��K�c�EI�Fn�����q;t��J(�t��N�ǭAO�$��JRO��'<^�!mXL����q�e���(�Q*�]�1��tC)�{QY[��y�M�/9�|*�t�QF����'��!fl�VK�zS�'�fE^�)(-�S*���q{H��`i��=�e&��֙I��l2q�zT5!���.l���@�	��޻n��&�O��1$�[z��=h|`̒��n�%�����7�,o�:V�ыB�
լA�`�aW=AZ�$���X���B���=`���F㚜Z	��T�i4�:vX'���!�R
����<;"�_�+n}�a��AE ��5��t?D��5��4'\��K3ɋ�M�a���y4O d���J��j��$nǌD�g�E��)��"�
.i��1��ޟ�Y(\����I�R����v�a�˞���x��TΥ&��`��
7w�g��-���y]h��1;�p���F���\K~���&(U&�<ᴤ����\���C�Hװ���4�	��d�Ȅ'����U���*�]�`j�
l������5��IhX��G/܄r�7>������Aoul�v�3��<�% � �:j�:����F5Kq)Bsc
zbڤ_���5ɗ� Ե0Y>��)�T�<P��gX��;��0K`2�]�����!��:��7A����`�,Y�A=���W"nC'53��,{�Ȓ�lD�F� Ib<OHA��tk����pܪ�wL����:�k����a4�K�`I�i]���v����E�'�Ze�@]�V9=�����dzB�H���g.�B��S��QU�+��Y9�9������Y�NR��t)=�C��
1�$�@6���/f�&hݼ� �̻C_�`mȏ�|�}�+��j
�d��&&~��V�]���]�/s6�S�f�<K�$s��Uڲ��sJ���0���C�P��̞J��|��2)�y u}s܀S����c�X܅G_}���O���y�<Q!��,-��?bgo��Y;������ []�gw����0�tĴ���Z�d�d�O�O��uQC/8�՛MN~���S����QW�X"�D�'��	ٵ.9���%��Xs�����/�Nw]�L��n����my���v�;dCF��C�M�1X�	%8�}�*&L��7�g �4�4�Yc�b�J�8�����^f&�vz��>�4�(��İ�|�	�@���Ƭ[�2�.�9��/�<��*n.���f��%Tg{8��I��.��D�c!�A�PRM��j�<�T�_�A��fG��U�*T�;l -�/-��*k��K9P�����^��j`*b��iv��IbAr*��y>aƘ�
5+� �sW��6W��	�7���^?�I/���}"ژ��.V|<:!+7.���r���^��Rk��j�02F?0���&��*�1�5�\&]]�+�|�' �\}^"\���C����
��oҚp"ꀆ`�K�(�7%O�a��l�����հ>64A��&��l��ee9q�G^���W��;�us?l�ɥ��1;-,S<���)���A���z���s:�f�1��?G� zd�O��6Ć4��zֽh���a0URVn6�И2�9��_��{)R,f�e=l�/���#����ل�����ʊvȂm��Ts�=Oz��B
���Ȑl�P�,���*��,DN*ZU5Q��>�:bXj�e��:O6O���
�|�J�6 L�,أ���GkϾZ�5�^\س��j�xi4x�aA>�T�zE��)6�&������%u��oy߽�ч������wF�K~�:���}
��[��D8��7��v/������U���L�t1�3�t�KT*�.\[C5�7�g��f�:�f�-@b�k�E`A�*�sd��o��%]J"���z(���Y��+0�w?��L}�7N�����x��GI�t��^�����Xmb���	qw�� 8-�9��1��j�����e�m��xUM&?2��1�⠋Xo���LPZ���C#o4Su�Ip�?u�~mg4�qb,..�9ΗKսi�XU��7⯢xU�ē�l`�3T계�����Z��~���i'�|P�T�+j׮�c	F��u��f�4�h0�X�eb���5����3�����4_��ӵ%�\bg\�� w=g�$�������TVR���8P"��䞂,�����c�83��qU��S���PC6�2<^8�{�6�Z-��y쿦ȋ�P���1+V/P�:�}�s�������,$��TA����Ocg��s\�=��� 6H�2�E{�)S$Em�D�k2�MeY=6�Ϩ��E=r������������	���
��	AG���HF>Ӵz�u^X[ȟ:k�.:aybl�voΖ�eB�E�_�z1�(�߾iB�O�@��QCq��V�L`���rD-E�b�r[�7�t���;�ۈ�^����?��K�n&:M��� HB�-�cқ;6^�6��J�̵x�����#�,�?��?gHy��'7�c|�>X�t��6�6Vr�.��9ӊ�Fvv�ˑ��L��6&����?��s�RJ7�H��J��b@�Lqf({��֨}Z�����{�@`Q�u�)��y(#A�n�����6��1�ы}cd	�!�	\]?�ǹ���'� -'��G�j�}DpM��P3ETw���x������^}�%$
J��7q�{6jQ/�b/'O��G��3֖X�꽟�����=A�j�b�! ~+�>t�
��=��l�@�`����Z��[�
3����=��4%��B>�C�C�#��Ҋc�S����э����l�*
�%��iUHu�3Z�#�7b�G�f��~��~1iA>���f"{9����V�톼o��5����>:�y)),LI����CG�֎���8�f1OO���m�&�7��G����	r���c�9�B�A�CО��w&|i񢒹ʹ��������ñ��i�闱P�d���P2h#���|�V,)��[3�����@a�2�)�������h���Â�<��zD(��D���̐H�F�X���Ԝy�T֠ՇprЎ�.��@:D��L���'g��mv����qanv��}�����
�F�^�fRi�d�\lxi1��P��+�| +�u�j��s��o��kQ��V�fR��Tjxim����f�q�&^�f� �B�JA�
�&�@��پ��ր�J��#"� (��"� �;�<��X` �؉0p�?d*@�&�LP��c�G�F1ϒ��N�i� ~���^J���n��:%�U��%o%��h�;x˔]:,g{�H �P!(�^��H
�?x���y�#%[�`�/��#�?aWuI�UY��w�͐�+BUg��TJ$,��I�ߌ�Ҋ>l�T5�C�V!\��<�z!�iw9U��/"�?�	��#��$��aK��1��4 }
�$g�۱g&�g2��B���V�"��)��j���W`X��`� ��c�$�t����I2��	�W���=�h+�41 ͹�S��B�v��A�!GeM?�s�Z�k�����Y�8�T�X=VB��9�d@�$�ԾLFυ\ycei*
^��Llbߴ�\�B/�a�5f�W�0ر�1dwi������/'�9����9��cn��%zR;M�΅���1o��i���K�XI�+25����6�Ae3V�g麕I��F;��Ѳ��J_����0�j�����5��ܺ�d;��j�`@k2	��`�֚)z����k�4�C̓T)�a30ǔT����~A�;ӵ���uϋ���Ș-|���:'{��]c7����*b����`?M*��c����9�j�w���]�B���=S�����VϱA�.4���?2�	�������2�GU��/�Y�D_g����K^7N�OO��'GQ��a��`c#��b������Z�g�l躚G�ٚeT�O?$H��f��<��GY���=����74�ۤ"��
��@��y�3Sה��q}5�[l5�K�6!j��=�����o�t��*���f;ZV9C��/���S
,�+ #�Lqc��F Y/أ�A�c̀�Z�У�n�ov�*W�El(�01�8��6� �;���l�
�ҋ*�uq��6�8Q�1a�ID��/���{c�$T7�'���0|���{@��D�0�䰉{��,�1pp�I*R�H�f�ş#�x9Y�nujab�)����6��ā{ c��_}	SR�b��Ճ ��}'�x%�H����y"���h��~��-�ZS�&�p!� !V��u�j��:�bK�*���y�7"U
5�D��}�F!��u��Z�*_mN�Jq�ke�\����|�Ċx��W����X���#	&��L�$w֩~<N��\���GL_�sZ���ǧ�s�*R�\��Ъ�e�*��:��"���Ֆt��0�;N�m!3I�j?@?v�P�H:~DK���"A���K���o�Am\���%u�j��\ދ��3�}��dq�W�U�a���X���rz~��c̠Z%�փ��i��pg�E�_0%�\p���X;ђ�.	ѱ!6�̄oɁ���~�F;0��{�D�"<�y;N�a�hF��#��}A���Ұ���r��`�ڞR���F���JǬ_�c?��'r���k�oh��`�K��델�}*�E�=��ᶨ1���|�*�iTn���$���x��#�m�������aǎ|��FH��$+�sQ3e�dХ�\���IѲ1"�?>��u)����Ĵ�6)/X 3�:���$΀򯻣����� ���8̫���N(�P��V��v����r�%�K[�m)K��b��������R �����_��������:.BmɎ��θ���i�-�y@��W�s!�7��ƀ��A5ȸݎ̙�ń�hb�4��9��4J�/,�y����-�y��z���kh��$
.��iZ�)�h�pX�5vNpV��G���x0[��7�tVj��D����/I�3�. �7H(}ͼ	,j����hx�q��OK}| #�\�l}��^�y�&G��?,�W�Sn��TU�g��	%B`���Z`��c���]|�1+C��3�8r�>iW�)=���a�?U��׉YT�r,�q1��č�k$�4�t�����ӣ���
o-�W+Q�ԉ����*C��z��&�7�qq�c���T`e�4,��zX�8������	<��\H}�7���d������0}U�&dE�����-FG	F�˩�����+�F��ؖ5:����	�����l^��NT  ��T�,cHzs��7Ե�40G�d_~�@��^�_�<��3S� �c�l D����ȹ����5om�G8x���4�� 6'��֒E��!�Ú�����Ϥ����r��'H�T�z�`5�D�?�#�S��%�U!�&%ww8�<����O������ѐDN�:��H3cd���|�&;�����C��v�Q	V��Dtl�qTd��bw�e]I���E�^�)�!Τ���.�b	��2�RҜm�r�~V���y�u��/�Ou�l,�;&|8���Ο5Rk��1tkΛ�p�*6@ƫ��y\L*��*i�%�;��������Mk��
͚dnï9im�(D4b���n[�9?W7.P��7��6��Nu% 0�G��WT'|
��p�#MW��*��X�4�BS񈉕�v:tF,���Tx#i���>�H_O��K��(�~U��g����##�a��l?�� e�g��u�y����)4�H�^��h������3NU; \��
��l��:y�D�`�����unlc���4��F�"�:Gխ��^[,��;L���(V�'1��W{_O��$���m��i�e��Z�m����Wߺ���j�L]�u+�Ꙩ��a��sZ&<��G8�6���E��?�>�;m���X�P��9�Jq��W����bH�y��HW��~�u���B^�M$I��L9LLUh�jQ������%�Z��@�/��&�[����=Su9(�A��D��q���v˩� R*��2�0`}"��V��n[w�b�i���躞�%&������<�����Ƒ��%:�OE�S�y_��|?G��{�(�ԦO¿�g�1�y��b�TIA sú�i�t\s�J�Ū¯�j�����?}C}��ǚ�}t�gÂO�un�4.M�% X�_����?�����u�2fD���LSg�8��\��.2���y�T����s�R����a����̌��/F�;3�7�Ѹ+{���#]�۶y�U!g�;�f��.�ѲK�@��[�0��H���^^>�%Ha�^��.�Y��r:�i�|b��t�ۮ�M��me��M�T�w5�����G�5��T���Ξ?���ݮ��n�9�"�}��[̑r�+c2�4��t������R�ǽUi)��&����?.�q+}����p��/l�LA��]��F��u�_k^��U�B��a��\�G{�xw���l�}�{���ZFj>j�VH�W8��P?�F������o���k9�Npg;+�ʉ�&o�Y~N�]pn|i���*�}���Q7/u����s���| �B���.�Y掏5����x55���_�x�� S|G܅ʶ�R14�ߣ�'�ܸ��۽��n��'�_����:�$��5u�(@H-7�OQϤ���[�z�7��GR/�80ʿ����qp�?ӈ;�g�����rz�P�ޖ����y2�K{�oVo]&������s��o�w�YQ�bԥhG�K���K1�܏'��s����^�-�"�4�.^�~̫}��Rw�u� �T =����b����|w�1�򫌻��[�:�)l�ޤ7^�.�����
曮:.֭m�g�5m(�� 1�Q��ۜ:�6�>#{}�n�I=ob/��/�'��Jo@SFn�-���5��Z�ٺ��J�K���6����>�ﻛ%�E�,�(��fA����Z��˨����v��J����MMmE�X]���˶{��+�e,�g���%Zl��Y�4�N�G����x_&ۗ��vU��q���y%_ga�����\��c��lO�w��Fk������k�E�?!��-�l��?���4Fybsrsrbcu�Ȉ70�Z3��]�r�5�������N�Q��\�<���V���ȵc�����۽�+��<��¡�ӦϙY<��F�O�F�[j�Q�.aC����w�����]��0F���l��X˕����������T�2�O ����Z�X�]�8�e�	������S��Y�0o�f�5~���U��ѻ�]�h�'Bi��z���N�N]~�M '�|ҼZZ�Σ��#�Tߡ[�s�(Y�n��7�X����yoB���������-��B��}�%���>V�\����$eki�h�V�s�me2B��ll�@���˅+pÆI�ip(��ϼ�����M7;�:��\�4)U�:xŊ7���Ds�m'^>ꢼo�b�iv|_�F��kE>NQ�4̾JܪܵIjj���Ճ��w�H�50�yom}��ysH慫�hIAK���緘ʂ�@�?��E����w57>��Ыv�E��(J�����%Gf�c_W�v��M�Ɲ��;�j��X�λ%*86�;9~�f1X�#��y�)]U��KnpI�R�|��� }�1�J��9u"�3��L�Ě��jl��$j
�����8�w�����8�G����MV�g'j	���r���&J��'&�h �o�J*jō��PK   Y�U���@Y�	 �
 /   images/8464ed5e-37c3-43b3-8b47-7240858568a5.png�wXSM�7�C�E:�	���һ�^,� �$�P��"
�A����E@@DAQCTPQA@P�����y�9�{������o֬Y{͚��d{d{`�oja
@� ���9>
;_|���)+(�֔� 9��C< (��ٿ<) ���PhJpM%U��b� WV�TU�U?�zI�}���[X�|>���y]C�w�f'M���&���'C��	
�Td�1�������`0������4
 ���;y�dCl9�o��2�d���D# ��B/ � �OP��	� -��U�T-)�w���@zG�ݗ��xoGLHh���
$3v�h<���s���	��B��g�Bp?J�����vD�q�n#kw�]�j��)��b5�?�f��� u�m�Bp?ʋ�+��C���B����B~G����"6>!a�"&�ƿ"`]�m����a�]3C#���h����O ?��/4À�3$���q!��!��0 �wtb@��."@�p�'�>�
���!�_-��ǎ��e��ю0�!�N�أ���K�#����YP|��/�\���8���CNp u2ć���8�Y��U���������3��g��/2��@�vu �	`�@~>wZ��Nڞ�%Ћ��ki�`�8�v��L;T�"���k�e'N�Sd'�$�Y���ޕl(z{�)���G�]ʥ��_����������Svd~��A?��{��''��O۱�w�(�w�i����%#��/�ws p���z`	U O ���� �Dp@��C�'�ܵ¿�?hd�d��%ï�{`p��JAV��C�֯Q!�"w�?"��jٻj8�j�;��&`Q�K���A����4���N����4>|h�_H�x��kT5q$g�ݡ�q&dh����!���A?'�]f2��b������PB�������bM����B�qB������a"B,��N�V?8ڟ�0���	G�>?-ż[x�d�u�od��G�!��v��俲3x����?�˺����WY<���������@C���kg��:�< ����פv󑛳��α�U݉�9 V�&�^�@8 oA�
������h��{a<����<�g'�����G�x������������������������������q'�x�� ab``��ĲgǞ={8ȷ=�YX��� VZP��P�@�
��B�_���~�������
J*jZ:z��! �g" ��@)()�h�i����`"+�R�Ne`�d	>���ȸTk(*��p�KY�p��x����"���u�q�ڤ�$Dm���R}���Щ/���WN�<�pxz����әﰄ��Fҳ�_��\}�O�/o�x��+@AjK��5��
�p6JP�`v*�����,(�yMNd9r��*���dh$T�A%J��M��B0o~��_k �[�� #t睬�PҠ�TöA\�������� q��l�����B�qx|cE�]fn�|ΰ�~6G�
�Bq:��u�I)+a�J2���cJ�S���\�����%q���2^�8:�8M�����!��1ux
�vn�g��\0����way��(��Y�f1�+Ц���^���}��/�si�����6
\8�?����!�ت���k[9߯���,���z�f$>h����*4�I��:���_��yl|��6���p����,�Jߝ�I�8=Ʉ"3z���[7y�^��o�����mjzX�#���A|�ڞ��m=kB�U�w���ݑ��n�4��2~�3.����~a�1;��}��C|�?�D�@��'AJ��~3��:���y���a���ߛKghl��l�ϼ`[ڲiy�j�3�cU�ʋ��-���]kW�揕�zW�Wd�!Ab��E߯��|�=�U�Ү8t�p#����b:}�f�M��6�w������#<ț{�9Lɳؐ�j��?�U�j�ћ�{"-�G�����b�r~�Vh��1/��}$x-�5���������}[�5��~��������[;h+N+\���͞�4�W��9og��j���I����:��[���B���;o��ӟ��%�������W�>T/=}��λo�qy����C�O���^c'��ﱊ�I7�;�7��?ϬE�r���\��ף/X���)5�V�z�C�����m��Z�D�>
a���Ϫ�91A��O��E��,����G-�v;b���������^�P���S^%7~����/�۾����<�ƄlP�hǎ��aj��=Nq!j!¤P���xCj�ɔ|�-v���J����m��|��[��Mi�۳�aE����D۲���Q����=�8�$�YT���n�J��==�S�5���h���~�^�tN"��0/4�����JQKJ�;�騿r�#�G�v�G܈������vJ�b삗l��2��k�e��Ů�x���1W�|Y �A'~q��!���Tu��7�xS���ҟ�ȋm�,[B����c��֗�4`c�}�ýᖷ����f����
�2׶��mX�b�^lf��T����v�獶���%wN�6��G5�Rj���,�����?(�iS��q��;��/ԝs�)��c�K�oU�9����~��ҾFB Z��m?m]я-Ͽ��
��y_��:`[u�G�h��cI���c[���U5�:�̀o㐳Ҁ��q?���k_�c�+,�/��ѭ��x�����w[���"���\c���T�x��>���/�a�R��<B���⍚�֜�����!w�?\WS�>eҿ'��������	�a�>?v�ho��JO^��?�KI�!�r�}��j��m�;ޚ��S�=_*�{L �|Br��<����&:[�:`[�p�cS1آm}_�T���sb��y�B�ܶ+U[�i��C�?������ﶾu˦�F��g�zT=\i��U�
=���٥��ӹ�㭤}RǏ���:��b'�e
=�iF:�}N���S��E��5A�V���亐��T��u>��ᥗ_�4�Y@Q�E�>/��6ϵ�Y���lV4no��\�>�6�e!>*�A��G�2���n'��=���D�\�9ɯ҂@�U�蕺6ԅg�/T�v��\��M��-ݩ?����z�2��6���YLq�u2����dQ˟��9�Y7����ݙ��B�ͭ|]k���4�����M����N�uI2X[߿��7��/7c_�Y�~�a.����B�_t�����Cφ�z^rŞjb^}4�X����~��ӆ�gP���g[|���k�>w�~]���mv�����!.�(ټ4P��<��N$yV%��$���%�+�!8\�p��%Z[ϴz�`�E��d�c�?ËԞß�,�^�pm��r��ۻ�d9�����;�\�fl���Iy��"��#Gqyѝ�����m � �����p�ٙ����M��{{�Mf~�]=>�[��#[A[U9�6�]/�O�P��:8k�l|bm������M���x�(��Aq�N�S7f�ږ�j�d�Yh�}{�s���ZS_�O�|[sg��X��gv$�� O�ll�~�U}2�y���\����r��a0���*�:�x������5�-�ꍯW���{u���>�F�K�.�|�g��|n��n�V�6�6��Hg&N�;vais��١ۀ�=�>�7�/�U��ul:�2|�S=[�hzޚ�w'�����&�u�k@l�6 �Z��xq���T�A��w��(�:{�Z���6@���ҽ���i]�T�=2�!>i���a��Ys��6��Hϋj���QF�,�V0�D��՚G���^6��^���o�'\���"Z�L����_��nhX��k��z����]�#�į�d�<B�7���6PW%�|��k����s�P\C���M�C��]ܘk[Ͽ?-��]3��=���k�ϧXIJ�\V;��r��ЬfN���3��IUu��P���ѫO��4�k���#{CR�i��=��rpx����S<���-aC��k>��=���3��uφ�1��e�n����k�4 �1N������zbU�jة���%�C��^����si�	��5?�r�Zq���~x0����^�XA�=Y6d�rC�b�A��/�~�lx�Tm�{N�>YR�~T=��fpd�?@L5G�Zͬ�f�Χ�����m���Zہ��?�<�A;=k���6Rs_ {�٬oi�Z�C��+V���|����h|�m�~�2WqU�&SQ��>�L�2v���9�8���@<;�ͳx,�k]�q��T}/���9������+�s��FR�m�fO���x����hC�7�{���k5��>��>{zᢼ�3��ƕ�4v����.)�ڥ����/iZ߽?hS�X���R皾�#�G��m����^߶�������&��2s�.�=��0��>ý�+�lة�â��Z�
+���e�=�tʱVMc�b�[Y�ZPEM��e�k�U�8Z��Õ�V�E����jǞ�y�n���{?�0�)�t�xq�e,i9D�������uvwMO	�	^(�ȋ�ذ�4Q�`�W~�ص��I�����n��I8��,W��U~��1��Ԑ�FGM�}��m�
�z7����:D�+՛͖u�/��.o��!��TNk�4-W�m�m�g���<�'y��x����N����+'�mᗋ���7�S��4G�̖#Jַ�u&�F�ƥ����;����3�5��n�6�&�+���*/>Sj�c�Y]�:�ڽ<Y;�ҵ�6�̷�<&w�mTH���5ɩ�Y!�����͕���4�Ӫ�C�I
U�З�Е����/7{W��.��;&����?���~(�?�������-�α�jy��[�iK[��h�����՘k~W�>D�x�8�X;/R)�]���ܶ��n(m���wH,�)�R/Q�x��W��#'[�ls.���6m�E�Rb���	jL>D8�<����\B��(����m 2{�|YH�$詨������6SlR��_��Ѐ�<�-8@�(��O��컟���R|�,�ҏ#�A|�s\�z�}҆�F�=�p�ƪ�T��N*������{�g5��5DvDfy�6T,1W?��r#������]ۏ8�X�P�##ZE׼un�7�>�<�1��ӓ�ן�Qz��!Gw�EwO��f���^^@��\��g����C�r�b��ևey�� �\-5-	�Y�V.������vXj���(	�(M���;�!���^�_�e��3�tx\$6���
�ke�d����4ɺR�i��߃-~V���b�ܷ��������	d�3` ����/v�/�C�����G��0����r���4S�zSi ��wmOr��D`���Bf��ҡ;s2�.�� &�h'��~���OfŎ�� ;�) ����~�/����B��g���&����	刁O�b�+�LĞ���Qo�gv�P�c����������:��:8Y����k�� 9Ȯ:?�;�)�FF0�g;��5�ő�� ������@����';6	 �Į�[��E?05��ș����ɶQ:�|@:͎cM	��M�-�0/�,bH��5Sd���%���������4�����i�O�L�^���w�32)v�C] 2��������H��-@`r[�{�������[��s]�C�������arY~бd;^��?���L���C&�t���V��G��"�b�� �T�O7 D�z���JW�R��RU��4��~��!3{������^0`���K��������&\	����9��ޱ��z�`��8����#��f�E�� �O���Taފ3��������Q�(Y��D�G�����$(��� ��� �)~`8뮴�w�����y�������������?�?~�����y�������������?�?~�����n�at�02�s�5��2���2�[aqx
 ą�an�0�~���8  Q� kGS�D���F������v}]C��v0�XQA� �ؑ=Sh�x�����À^�dLA�.q@A�M�>�Xn�g�1:�1Y� t ����LX(�<)�
�	aXL8��A,�1�`2G I����b!�/��@�Hpr0�> �e��{��C0;G͍�A�;GaR(i\SSf�	�����!Q�Hf�B�"`��;��l[hd5����<B�������0��v}����q����;>�e �Xm���� M� ���o��E `�q���p�ۋoHH���bxx��R �W��������~�f�{�F�
�%��AH&��F�������s�xc��leX�X�84����_U��2���n���-��S`� �s� %; =xL���7+:���\������oΝS��oD��ik���	�
%������f��Q@
��:��&�~�p܁� 
�Dǁ�,���b�
P\�&�p =�c�)0
L 3�G`�
�C ����Cd!�Db��8@�!G >$9	9Ʉ�C.A* ��f�}H�	�d2Y��Q@))8(($()4((,)�(Q�PS���H�ȥ�LQM�Hq����)��G�( e�rA���P������1�$h�2�:�6�:��~��RRS�S�(�)�)�)�)Q���1�ɔ��W))RQNR.PnQ1Q�S�RiQYP�Q�P�S%P�P�Q5P=�zJ5C������Z�Z�ڜڝڏ�u2uu�=�'�S�+444<4�4:4�4H���<�j�6�A����B�ZSZZ�	��J�V�A�w��t,t�tZt�th�H�4�+t���f���Y�%�u�������_�D?F����A�A����ǐ�p���a�a���Q�ш� c(c*c9�=��_���$���<�B�R�*�0�f���}���=�=�{
�4��3�L�,�l�|��(ss=� �':	#$KKK3�s�VvV8�-k k2k%k�{66	664[<[	��)v(�(�;��$��G�3��~g9�q�s,p�q�p�pFpp����rIpYpp�q�q=�Z�+��`/fo���{�~������p'q�p?�^�����d�4�����������6�/����%?���1��^�A3� �<������[g�؅t��B�BmB`�0X ,�� �/l.*|I�_x]DR�Y�H��+QzQQo�l�v�1!1k�(�*���t�����;ĿIHJ�J��h�x/�-i!yT�JrL�IJO*X�԰4�����t��c
U_��Y
Y5Y�l��9*9M9��e�����a�U�
\
V
'���=3;��T���(������'��K
Q�VfR6U�U����"��Q��2�ʮj�zZ�]uSM]��v]mV]L��z��s;�d�NM*MC�X�;��ZjZ!ZuZ�����+���܇�weߔ��R�΄.L���E�	=a=��e�7���h�2�w�~��J���oFZF�F����f�I��&l&�&�&�MEL}L�L�T͎��3�2�4�0n!`����Xد�?z�CKFKG�|�7V2V���������l�mp6M����m��+;I�`�{j{;���p�(�GvGO�JǯN�NiN��RΡ��.�.]*\���f�N�)�E����c�oy�x�x�y�09p���AՃ	��<q��0���w=�=���G����<���E^F�xYxz-��P�Q���l�,F��y�����G�'�g�W�7�����]�3�+���o�_��PHx$�ǆ��=��#�O�d��&����/,	eD��V����
=:�V�=�%�>�5�)������c��P�ڣ���GMFD_���xŴǊ����ę�]=N��x�	��'�O���/?u��TUB���ڧ��P����OTN�K�JB'u�U:�sv#�ܝO�M�N�N�OSK��N��K���q5�5�h�T�uVc6,;){��繮������C�O�Z����K�����Z`XPS�_�X��]4xA���b���k�G.�]j�,q9���$����+��e�eg�6�q�W�>�P����L���
���>X����[��_��9{�z�C��gu�u����o��,l`oHj�4F6.4�6M�r���ys�m��-
-�w���弛�J�ߺ�v�m�^нO�}�O�{��>p{0���a�#�G�$S҃���N��;]Z]���M=j=����}�}�j����k>��dߓ�A���C�C�a�ឧ6O�<s~6�������/_��\��Kz��*�5������5jw'�'{�8��BM}�&No�Ŀez��N�]�{��;����?�0�1�����9ֹ�y�����?�.�-�,�����|)_VYn_�[y�5������<߯�j�v����[ߠ��ݔ޼�e�5����=�l�c�#* �aP�@�d�"\AIا.��1!0/��#�M�E눸�Z+Ya|��G	ǣ6N���(M���.l_�VD`P &	���"tDv�k��LV����잣p��MLUAMWQ��k*�ՔU45���*4�4���p5-%�g�A|��`l��]`LG䏵i����.�5���<�!O�ą #�qDџ��u ��C_9���興�,B`�/���V?��������9~q�<?����J��+@]���{mqCL�B�{n"�'c�"�dFaL�0�џ�Ѩ_y�B	;�D�1�@����*Hˈ�A�`��KG�|�A^IU�p�y��&<�	��Y�����\�x4�;�_E�8T#������l_hd�d�A�C�"lB�0�',v��08���#�XE���SM���WD(�)k�k�=�;�����Y�݌�H�/y�	
@�[���Vد��E.ٮ������Za|��H;'#c���S5U#8BC����P�HE	a�a�l�l��0����{�焠�AC*�I�02�#ཱ`¿low���Z��
%7㟽�Gaѿ�����R��,���Ǩ�x�#�j(yUo/e\ISYC�41�#�DUG�(`AIJ���*���p����
R	!���T�W� ��(4�ϟ�w���S+uuC�����������������2��D��HUICUC�Fiy�	�H�n�@�F�/�C1v��c�`[��1�8b�� ,l��i!Q�5HD�a�"?��Soe��R%��)����&樓T��PAb��?��bpo�Jp-��ϖ��F�{��#	���a_�͉�E�|ȍKQD�]���r������?.����R�{M*�m2�Ig���S�.��O�'��	��������1.-�����(`@��@A^;��7� ���O��8�_��vC!�?�/?�ȿР�}4 ���T4�t�� �~�Yf(���PP����eV6jv�VX��NΉ0��W6D�6r8N�-��q�>���#aQ�	u�v�d�eP� ��Q�_o�������҃�v;'����!�4T4���.������]��Cn`�)�@�q�XS�T{���ד�EqcG��[B�x�r;���	��_��݇�T	��^~بJ�8�CR7�kzA�=O.����C<2W�,�m�m��ռ"��MM�r�Hȃ�ʢ�Wm3ɔ|��H��:��(c����x�q�i!m�ﺹ�dM�m�>�v]s禞�����f�*���lD�� �gV������HM���H����Yb����%u��
����e)_&�jA����Nnaq���r��a0�lV�����L��z~f?a�����J\��sa�
�����jЫ�)�p�l�i��ߗI����)ߞ<���O��=�2�:ŠnC��|�6 �<e��[�z�"�A#q�𞫱E���~u$c6�6�^���VUV9�+����RT_�U3����ņ/��)q���~a���f08E�[�6�G���ɥ|?�i��L��.�>���>�Z�z�,�pb�3�i����>��{�Z
s�7U�t����L�`!~�  u���(��QT�~7��/k=����H6a,�����2���lz#����<yn���}R��o"�e[p����GQy!��o�����'r�X�d�h�;;DR�-~_����j?��(�u�}��	�1����s'���2ɲ{�h�4�i���3�7�/*G��H{\�0�q"���2��x$������ĉ<C�f�t��� R�m�ͻG7���8���O�3B��"��H�.z�+��9�ؗR����}QQ�B��Y�;�@���7�[�	�O�o�j�[�&M�>G�$s�������~���i�z����OU$�Ι/yP���U5>�z�ž-�^3رq�(JB��*�U'���W����E){q#x<F�8���U}J�G�T�����DB�~N���B~�-��ځ_f����|�e�n���c�E�S�2n����$9S��JFeh���~�*y"PY�X�ݻ*�e ��k�(C��*���\Ax]�xT�Q:�VJ����+��Nn��&ߺٍ.)�$�V��$I��{}�Pr����m`j�;��ÇF�����i�-��U�IvP��	{�^FÓ������?J�{z���T�	�V��_��l�d�{P�b
B�i�pt��Oښ�ҥpa8TW��SZ�I�^���HnD�����O�Χ��ߤ܊n�ԍ��g`�2�P���Y��3D�W�{p�C�1�V��G�� �*�kK��ke���,)E�Ä�D'��>����J�K�;��5�)%6&��v���]�;Z.t��2��k��ؓT0$t�J��S��R3����,DR0��&�v�&%�e��QO�⸱KI)�O676pj`נw��2�hU:�-f"@��Zԝb��)���9�-�	���pk��i�'���ȧ�m1�>�;��{Wb�*8�M^8_���׀W�A����ɿOF���vnK*���k��`�m�~�(����W�����@=�k�L2�
��͵�2fX��U������3���-Xڜ�6��fiV�r*�ׯ�X��X�	{uu�D{3��l�����¸�e[1NE���K3��6��gG�U�-�r?�!m�t�`|TU����wU�k�#h����U�4+��g����,+��B�U�iB�0��_Q^.s\K�F����*χ�Y�8��au1�ܵ��i-UPqƴ�� "�Qp<�*�D~N:
���:�z�N/�1Qv�)e~U�P���u�����[�d'%s����m@0�C.k�:�J`Oߡפ�L�N��E���LG�oP����չ$�t�T�\=����hj)��/5%�ND�.a��|��6��bC�J�k����1�����+�e�UÜSq�N�+S���V��aվ����"{W����3�T1�^�p����z����X��c�=��	�A�V�n��P�l`(�<�[���M�j��Rߋ���pU#�����S1�[��[R�2�E-_�Y�`�[�l�[x���H�T�����-J/r�5>�� 6�4ح�}ɕ�Q�2�t��{V=�]�f]���yl��=�b�Ω,	��`V���!���Ϟ��'��xf��v&�_V�J"��ULeޑ ����n��Ӑ>��`:�hK����&9��-AuM�	��`�ncZ��
�h=��gf���g�\T�Yx3O\�ڭ��~�~�<0��Lb�Ⱦp�s���l��c��o��Rm�c��������h�n��]2m���1��{�`Vi�;��H<A��{K�o^����5��8�~�'�Rz�?��a*����p�\,0�+�ר������+�P�ż=����i���}��=��{�Te	���⯯S�UG���h?���{_{E��k�;�N�,.�#�{��·����ȩg�E�)�V���5�S8����׹^�����vuH�`4˛���xW����
.#LnƵ�W�ɭ�l�~�i.��z���q�E��}}`�I5�����紵�rSy��;MS#�z����Y��IVw>ǰϑNEM?^�˾0�<�<� U�8Vf]S��C�Q�g��z���# ��g�G7I�n����w�>�wnx�<��:�\9/�ª��Ƿ�R���QV&#�a �DMܯ�ԫ
����y$��	;��R����m M�97���3�}y*�O�E�c�GQ{9Պ��;'��������;��v�Pҵ��X|QZ�R�;>'2�/^�5�F[y���}x�d�f��XC1�U�^���/e��QX?g�*����V�Tm�3B�r�}3־�*��	6w���0�ZN����7�=��9>y�[=p�$�F�K���E�/���p�߅��ylze_9}�*����HY�*)���?�d4o��.�Te�Zڊ��P;��wg_{��iJ�O(i(Ny0�B���b���D8��ȯ��w�����l{p�n�(�ߧmr|$EB�	&���\.P��(����[�P�]�������ΫU�{�����p1p����L�����ʩ3�<YY�B7�e������m]*�f:����)��wwם���ԟh��{�C<�"�*������:�/��ձ:��;�`�{�*�~_�C_����}�5iѴfSV�i��{v�O���f�/��މ�Ku,��G��f&�{RĜ.S���ydH����f�L�/^U>�t�r�>�W��.o/41)b~��pEm
.6Lo*��:�h��>���VqXO�P}��x,�u��\W����H���칔�*��g6��<߽�vy��Ւ�8�ɳY��A��>�
��W�*]�'9_-�Q,m__/n0ET+V d�0�����A�I`~�pl���{*.��ʉ��L��V�qqmTM|�4g�$r�j磎����y9���|U�5����c��\ҥ33��#�*�=ﱺbfY働`�3��wst�w��쬍J|v��0��E.�}���8��2J��qӜ�z�ư n��R�¶LI3b��%��8����rii�R����9�z�iu���N�J�H��,�F�ed�C��ߖ��8rj��R�\���;���g�V�<�Pێ%8���*�?\��|���1f+/ڱS=��l�.E����9%���W��E�m_���QýN��wو��ş#"�a]��-袟u䓹vb��@BՖ�6��o�f��M>uCd
u��3��hŌq� �Q0I�^Z�Hm�U0�/u��T�Q�´?�nc����S�>�u�5[�N�Vә��%cc�#%�[#��~�W�fd\*�"9��]}���E�������H,�p�����O�^&^�&�
�2�0�b�tp��L
c�|��y!j�<�qX�i�'���up(�gP3r�I�����"Cj�4\�j��~�b�7�b����0+b������D#�����T�B9��:��ۮ
��B����O\|
�BOsȷ,~�[켱��\$AK�$U���}�i�1�[�F=�+GQ����~*�-"��gb�$.��3�7�S�Zo-Iw��R�-mі� �V�d��
h�Wy�(87IG�wy����ܕ�f$j瘲�:�Ll��IH��m��&�m�C�Z���oY���ْh`���QmW�d�ˢi]�T՛���^�<<�8O�s�z+����ʑ5p����#T�l��LH$P-rqi���4�<AA��˃.�w�]�J��`��3Ly�Nɜfu$�1�_�Q��y\��2�uqKj�טZ����jp�:�I�9�YY�j����a��cK8�)�q�$����ߣ�pO���QF�XDl����rG�6���8�!�~:�۪(��10��;�n�s��Su�=�#���g�%���<�0�2m�Vy��P��:�s-���:3�_��.�}�}���ѩ0��G��)A9n�F�"�4�T�u���^n'xb  ~6Ydj��ljV�����)���8�ia�^FB����՝H�^�G��{�����_���c��ƅh& ��:�u��R]Yr�m����L���4��Weo��!pmڐ�~��/�|Ȃ,*~��a�G
�i���	�����\v<{^Zd��m�ZN�~�'�Tu�U�ǎ6��3����}����ゕUl� S-�-����,=��d�S�x:�����ŷ/��J_$5#Y�;B�,��E��{��*��M��
Pz�G[cYO�=it�V��ǜoU�s=�賽+*�2��	go?b�x�z���d3��%lo|̝�]�~��i��&�T:���g�K�� w�k97����	Ϝ�+_�z�rZ���Ū�?)r�C߭CgF�ƻD��_ �yd][|F��c��1��!��]C
�Uz���	�^�<����^]�Uވ[���o�����ˤ[�\�a�d��G0<jlfh���mRn�ټ��8�\8r�$�3um q�GN��*-�{xA��K���=C�Õ&ot�n��=%	�m�/����+��iSo��k���P��
>�N��b�s�446˄��e8��<	�Ն���2:���U��}�nf��gc{���%ڭE���W�Ǩ��o"x^�M��E��){��\�n-���b{x���Q:��\�^7�,���|�K<��猬�w~�wWǼ����u��hږ	�Bgҝ/j�d�B�g��~�i�L�)�4�t�U�r���="��JD&c$���\kH+��=,�����J���CG�ē�чg��Y��O}C6��jW��:sG>�7�('�t|5(���'�q|M�M�;�Z�[�i�q����I�~w�{ǻ�X�bt���з���������߹�Y�ݠђW;}1U8�nD�
�EKӛ��>��\��\���P�����
�����r��l����$E��~Ǹ"������k�7/�,�C֎!���<�S���y:K��g���)S��\�,�"0�	\�͜�6��^|����ʡ�R������;���ĵ���"/���k٢Zb;����KL��Ov���5�Z������Od<y�Q��~����=}�l�{�l��ÎK�]�J�m�9�-y��%f)/��G��L�ns
�f�m��7��i`��;�P�s�5�eQ[�O ��_��j� ,L`:��A�5W�n���S'Ա� [�lrn��yN���U������I���K&�X��/��fק��n\rZ���Xj^����p��-�"�R��)����a����s���f�r�?��=�u�� M]3�ɉVR��{|*ї���Vf��-�:�
E_ݩb��׹]�QJ$��	eYQ�s��r7�_��}��u�bp�&�*�w|��O�ɤ��5����<�b������nh��o�-��U�k`�Pp�xȺ�ނ9�Q�	鄟>�%w뭻�ė͓���f*�G��o�N}�����1G�5������szL�����.�9#o}�;e���]q��|T�A��ϙ�{�E�2}�����	�O.��f}�����=�K%��d�Xa�j�/"n�l��T.�����2*��Ԥ�otH�k|ϥ8�OL�~�)��֧=Ӄ�j�*��\�*�:��.��|��;H%�1��ߜ6�����Ą��7v�V ��dF^C�n&�k����D��XhB����|]:Qpe"��O�����.~���fN��*ކf5v\���1�o5��(g�	�DN>�:�:��=�y��e�3rR��[���Nj/�x[J���R��칦s�r������`�B�=vG�2�4��(A:u��=ͩ)�iot+��	xڒt�ԩ$����|�]�I_n����L�7�I7���%E<�ZB�Ú�]V���+{T�eyj�|��Q����;�l�eC��dov���+���'�
�1L��\(S���W��1�/�o�Y��L��E4����6��ڰLڈ�A������{���"W�F�𤽬A4���~ZA��F�xM��/~�<U�+PV�!��|ʳ�>�œh_�L��R��I&U�׿X��r�q(!�}?i툵B��R���cI��uS�Pɀ�>��R;��B�J�)_Q�/5"�ڟ��s�x��c	��^Φߟ.����x��n�D������U��i$����b=Q���1:n� �̙�zn�����.�����K��p�Jir����H>�a�R{�<���t;w�KOa�S�c�D�����3�S-�^S[���^��ŧyޏ��ӟ��8�����E��hBr:�KM�K��Ha��̒E�����j��=8X�7��e̡�$  �W��_6�;�IgG�7[�~���xPy��J��g�t>T�U����@o1�.�x#�/���&Of�LL˞�b_�y�Cܸ<�:��LR�pcN˺�}��8�I��R���e�R)[lO@�Wg��n�.D8��� �Yo�}g�;3r:_]WoO�h|�{�=�ǂ����'��X��Δ�Cj%���o
��skW��u���KG3���C0v^r΃�a��9�!�I�
�ݯ��H��(�k�˗U������넏���Ӆ�1����唖^Ͽ_�uG�LDr�{�{�T�����o�^֥��������{3 *�7�ߕ b}B��$ӆ�Z��p
�ixhz�d�s�yV�ɕ�U�%�L�`���;ܒ=Dw�K�3�<q��3����CCG�h�x�
F��-B}�9b9E%,O��	ǳ��m��"�]F�Y�dOL�	fU��|dFi�ǲ7�97g�Y�\h���zA蠏���'G�y�U,��.����x�������3�l&��IO5�S?��L��0o9�!o��)7�f�b���c�Ϻg��9Ԓi�ά��	����%�f���Uy����%��3�>�8L�_���#Ώ0���䷼X�0db��iޞg������'x,��{� n8�{�νTg�<�7��K�Y|�rg�s�x�[�r%�upRI���羱� �勎	��
���e��i���!n�j�V�3÷��[,eD�չ���/,��:�8fV��R�{����U����K'n�ѓa2�@��$�M��%���f���xt�<�P�����7�?��>��8�X�w�\�ț~�s��S:���b'�O}08�JS�9�^���
Θ���#����RpϢ�a��g�&n�:�t���8�DS��gߪT�UH��f]�����B����B�Ӟ��Hj��K�M�ƚ���<6R}y��̾��88�����F�at��т�t�[@�� 9���=�t�t�ԊzP�6�c� �?��������}]���ϛ�w�ɂ����r���X��I�TaJ<t����Lb������_ �\.d����4�}��ᗣ"��s��%$�nK%���
�Ì��J���K�J������Ϥ�kho����_]k# `_��!�P���-\��?�\-����5�/�ZID��n3�W�n������z�����5��S���Zfc�#��f�iZQ�d�������[�#��؞��	!���U ���9�v������oڋ?�:�`F�p�;4v�vuE�@[(Ļ���ѥd�:�K&��'ɉx�y���N�Qk܊_f�������h�-���@[��߿Tl&��t�q��Ƭ�H��U9؏���MՖ�;��^�.�K��]�yf�M�"�l�fpX-%�d�Q��Gm��x�G�l�����ջpָ/��%��.nXu���?�}o�]H��o�V����?�����K��sg�ɜ�A���v�hy:M��J~$���ٮ�P�+���-ǷSH:_yE3~.!�
���Իá�r���ǁf:�de� ��RZB9��\6�&��?(�ۮ��w�(vgM�k5,vg�C�#�Q��\إ|�&Ep�`=,��~.�<�(��+S����
�����l]&62]ϭ�?�z���A�6�1��x�$!\�k���d�����=���J�g�S�K��fF�J:OJ���c����{�42�M��/~�D��pS�N��T�z���_ n�����D�s�[���Œ�CL̓A�;���丟���{��VN��c�M���I��/�������V�����\�`H�eT�k���ǎCwy�77)�s�?�]o03�뱶͐��
.�Wz$�签q�e�K����NCܓ83�X��?4u�Z���B������"ԧ�ui�p�L!��M_�f�WR}7H�/��Ǘ5%`������1��Q?<n$|��Se�;�\��%C]K��*]6�2����"&uk�S_�R���=}э,�����SO������5��WKŵ,�EUr��s[�1���s�P��%b�[v���T��5�(�Q-6��M�����йپ��e�["U��N�*�
��b���)ς>��Z�����?�<�v����v�e2��{���4������V�(��6�׸:9�Ul �:���r9�j��e3�4��W�5��(�lc�Iˑ�z���~����_H2�܀�Q-��U���"]A^�A�sæ3�d���.\�����+�oXS:S3�������Y���L]��-�}�Y7��sBxK7m���6q��3����2t��!o1�~:gVP�_�)A����ra��'������1س{��F�o�q	�<�E��4�L-��~�zf&�N�;*;���:�{	,��R�[uEւ�����]N ���u��Tl�����Ky�!D}j�wvw
��r��0��U�BŞ�f!~��Yئ�wu����.:��5)?���GW�ߪ0���עs��/��58�*ҍ3�ؚ��rߟ��S�:����?̄;1u+�֧���YK4;�?{��C�(�F&>�2Zw��9��3�s�B�a�ؚRD��Ӌ�)mj)��&�%�
�4�?����)�{�Ð�{��kNa/K��K9MGk���G�e@��S�h�2Q h�
%�j~�Z�.!,�b{N��r�����}Ў	�%Pg�����U�Tzr���5�a{�Г\Tx�3��^k�$�d`C���w��WJ02��0�n%?PY����h�9-�Y[c������Z�vA�Y�)"�X�;I��_�Q�:�\ CTRC�A�m�m.��M�;K�Me��[�e��N���F�Rՙ1��K��X_9p�~%�T���;��y(�ȕ��7eć��Vw�=ړ�Q����w�H�gԮa[��ҞR*�Ҏ��.Ђm��zp����}B�A g֙�����,XE�K�);&s���y|O��q,��(p�Y�,�qâ((��+H��x�+0���s�g���+�M[�u�Xa�o^nX{4�x���X?Ce�9;��^\?R��(��,�"��6]���&vo��iK�1œ�D���	h	��M��Oz��(�����_B�?�����!F8�9i���X�˰x+!�!g�#0����<����]�EA٤J:_~�6fTb"�?[�}���2�Gx��� pFuk�۪o�d@oh�����:��c����ec���x�pkB���䮥X��+��[|p�]?���M�@�2�
�ӇV�#J�������==5
z���UO����{|�S"hU*��;�\�y�QG�jL9LG�bdi����sБ%�~>�4�5.3�ƫ��.�ﮆ�f���(�d�t�XCZſ����{p��W�H`��
TMbQ����v*D��c��l��~ݕA��	�w��e��%ּU�6>i_cxx�~�������Y U�T�u�F޾�n��w0iep��p�_\EX�07^�qG����:�b`�;��5��O|NU\�SeW��#��{G@//�:�CP��"�}Ba&ӄ����|���ؿ�����SxQsV-%�.d������3���]�d,=�](YѰ{9R<�4�Ĩ�5ؿX���j��{��[���\�1����0����>�}�������?�f���	�81���>pR�F�R���*`�ʕ���@3��B!�./�ק����8�JMv�fwd���OUͮ��g��=uN&��=��������[�n��S�!��N��Ral���WyGк�KԄ���8�]x:�~�.�y���.#7�u��}�$���"G:�*��d���ٖ��ᶤ^΅�3q@[�����k�K��[�� �?hZV�̢�B��P�"y^����v�
sZ�����s,�L�J��_%�("�*�iYyd�jҩ��Ġr�\�n���=cn|�ѝwP�H���mt�G���4���v���y��r:ː�P���/������C|j�� K�5֙;Q;���ްjh���O��Q[���^�*ԝ^/K[�/��y,l�؞�=��}[�EB�̀p)�A_��8�����j�%
,	BE��V�I�Ʀ��k�W|��c~�sE�K��n8;�8qKD_�NY=̈́�ﶔ����I�H.Ĩ�>p=�Q�1#�y�25��Y��0
O�^�b6c*I��L�'���fH��b�*�RyaȨ<��{��{O�(:�V�6^u�$]-�<B��ȩ�"�/H������?ms����]�q�r��JC�A2ۼ��Kb�թ���+��@��
��z�b�=GY�v��E��f�ywz��*���A�c���� ���J�3|�t�
��=�~Ѵᾯ����Á�`7N�u� �V��4���y�Bu�0]��1,�(��W+��[ �������4?}����w$t@Z�e=ԃ�
vv.Q�� ����̪ �<~�a�'g@�,���nݐ���L��F�T5�m���]@�C�!Ⱦ�̯�Y���p[�yt�G
����:��{L�[�5TN�%����"sה$T�7�7\eP���M�iv�,�6��u
�o�M�CZʟ��!����q��_v~<�_�;b��4o�qʧ��Gp&�f3�@��;���-�$�,r�S��I�-�\�Ĺ���:+�2����C��K�����ӥ%�gb��)"��C��C^w�Q�ۢ����y5�a/w�X�`@l�Q��\i���3ENy��>m�����Y�y�<��#%�}�谛p���۫@��(��6s��e|�d�DGu�5�>�tnI:)6YMxߣ*�y�rxv���$�/$�ؒ�v��x��d����d�M���%1q=�bh���,��H�%�rr�w���ΫRh�H"߭�w-�lVח>���ߴ��~=�D���������t���p���
��6
��� u�����޸��]4*�⻄�Vp�W���d�p�&��ecC�܆��TGK���g��W��()��#Dԑ�еmU�T��� p�6���i���px��*��;iY2' �{�u+n`SPce��fl� �N]�N{�h��qݻ�̤��]����e��:�uش��U�u��0�9�������L���Q�}H-��lwj��T�aeٯ{�:|xa�7��R�Ӝ7�#��M7�n��z�xy��vo?:7� Y��u���)����]�N�&�_ �"R�@~c���#J��)|񵾺����!AUŎ��c��خΒ)���NM3�kC翈�5���K+�c?�g���6�u��%�����r��,�I��^�'c���^��9G}o���m��X7�����׾.U�h.�\��]���	��f5�w6��#�{{�kw�,%�;@K��$�ؒa��J�]�y� �y�Ț�`r�e%a��|�kCs������Mo<���|'���MX,s4t����/c��LkQ�Z8fX��/@3a������PGkC��4�n�z{�|wK�2|������5��z���ƺ���+J��pI�����ućew�����ğ �=Gre�gO 10x����6�v���Ǭ�n3rP,T�C�2;]嚯�ۙ}#W�/�[�s7�\{�б��W�M�ȩ�(g��R2�j�u�Jk��*T�����f6GpMӋ��^�tk,c���A��~cª+�?�s�uu�x6���^�iM#�%2�`o��Y4�_c>s]��p���7�K�W����`#n�zgҥ\ٍ���2��y!L�ڑ���~/��@�$�8��0��vt�����_:���4�\���m���)��c�yN�B[e���Ap���|3o6�3����������p5�G������N�t�X��@wb^/2��%��|#�BlN�[��a��v.u��#�{PU�Wߧ��bO�W��L��Ĉ<�S[s�tԼ�n � �V�����S���p��
_��1�\8��[���*83���� p��W+���j�e5N�̢�͒۟���d������\��(�.~����s�����b�],�W�+˔\ ��	�h�x?�V��ZkV�}�K��FI4���	�`�0?w�e�%��P��
��;���+�^l6��x� ���?���h�ׇ}J�JnᠼZH�m��6�m���W��D(F��ٻ(��$�3��G�}�	_7��ڒ�J��Y����0P{O�BV��;��E�~_�w�c;�����N�Ā��Ј«P�w/#��,�w�+�]8�`;¹����i��_N��guP�r9�5m���� �{�FK�2��^Z%x\O��f��h�_���� ��[b`�븯��+Mr6Hg�8l��*�A1ڏ� �#5�N#��h�����_@��;4c��k���� y�D�Vx��T�wK��DoP��G�$�Sy�@��KWR�4(�F�5�0b�z�����YR6����S��<	�R����|'ؓ�H�|Q�'�0(��&��������>_�͍�oa�!+5gd@�W
���yS��!��S��<��L����g�ݟxB$}�;s+�׼���m��H�2��4�A�ߠ�C!�uB����L�%y���e��1[(t#�>+_!�Y��ƭ9��d�U�uȷIZ�H��9���{��K�I>�`ǸC�L'�2��|Ai�h��j�*	f)���Y�c0����R큠Ivx��W�Oo2�����+P�C����S�EQ�c�U��Kb�4�Q�\!V_�^��~W ����E�hb&{g��P��wg5� Wk�A��Aފ���5.���fa�	��j��I�=�~�"Mߦ<�2������cŷ9�G�H��I[�Z�ވD��?��}	��/T��4�;j��H�hu�)>�q6 ߆5V�#�Kd�hg�_�[3�w����K�����%����)�,5���'N<�}'��9�ce�:vR�,!���L��wf�#����[O�`͒�t	�	q��z�Mf�]�Չѽ�^9h��{\SW C,����|�lËl���Z�C����9�� ��s�?u`\F4��L�n#cS#%.��}}:,����+��I�l}"����d:��D��+߯�� ��k�z��A�}$�
Н\�5v��w:~^d>�z�y�4�gr1ʺ�p�,�05Y��B��^�S��x�-q>��qae8��;
�=yf�?�q�b�Z�d�00��B��oШ}_�Z��yl��k����X=x�����4�l�=&�!Y�����b��m�z�N2�v[�H�)85ɛ�-%�}��eo<oa��`-Q�7O]�(���@O��b��#\o�g��[��4�G[)��J���s��6:�5���`Nm�]댩춮j��jӾ�].(�e��������$�w������4R�F�uT�mnӛ'��6�Ņ�J{:b2ɏH2}��@ե�R�A�@q�c�F��[ل�۬���4��j?�]'�H�6z�����)�zUT\�3bGtO�ח�r�Č�x��Ԅ�R�z������G޾����sۛhS�d(	7b�x}7n�Vd��1٧�)��>C���^bV�-��L�6�מA�q�\n֛��g�Y��d^�B�Q3s��Ɠ�������TJ
�� {�OӸ�?YG����LM�X�������6�O
9:[�2�'�5}�o�L���)n��m�B,���&x��ė�~���D(�L���o��WZ�}M�I� &��3_��ènm�X�*��6�$.r�/���R.�%K'M�>"�c��TE��R�
JF��?�{fe\|�P�Gaod1֞^� 7K�P�h7�`[��}"��� ����3���Kb�]��j��� �> �{������C�h�|��F�����lN�s�B�������,:��d��J�7��>ϩ���H��Ɇ���w9���q� M0e�,�nu_ۍ���K���&�/�U7*}�):Z]�X��n��1���%������Y����h��d�5�!�MF�,�RBN��i�
�����
�ڸW�i���ˣ�?s!��Մ�-o��n1l��[8�	#
�w6(r��H�R��41���tMa�2?p�'m����rI��@�{��N���K~Dq17�!U`����w��}1�b��IB�϶O�A����I�~1�Ր{ݻ�5�H'�k�I"��t8v{�?�jj#~�pxB�)$p+\s�}�?x|�s�6�^�����%�~�,�D@��h���:�yM���g�ʺ�E�*����!��#x���2#��P�x�t�@�Mz����o'���� ��`N&τΌ)�=�U{�v�q���xK��w�?�@�Rw6���0��5���N�m5i��ۭx\խ��%0��Ii��	N��k�S��oߍ�iUDM���R@�r�B����j�0d�H��!b��\\H��P�Tt�2q䳃K�N+�}ѹ�;���mgu�E�V~h�y�0�e��LaI}s4Ǽ���CR�$�����N�c�\���:��3$E�$VF�BI?U�X��e��
�s�\M�( �]����AU+8�H�c!__�`ٟ1�igu7�L�@�7��;ݕv[x�V�ڹ�\w͊�M��
)��[{���������?v˶�ʾ��:"��ڃ�/͡�%M���H_����V�Cۼl�b37_m!U��&�h%���+;DV��
��{�1%�[΃Ʃ5��d�qx���R<�mfgm�Iߡ��TV�,�+I�������Ym�˯�>�@H�^��Jm��|�R�W���ZA��SC�\�d(mɞYr8�#k�+A���	ѭ4�^2��2�/U��ܳ@jd�ڀ�ؕ8��>�_y'�N؃U���X�5�`l�ۼ�Ѓk֪���a��ə~ۜ�<��^:��N�9F(:!�!J&��o��J����T���Y������VԔX"��{�'�_1X��8���(�?.[�����(�u�Kz���#s�@���k��ceޛ��U�B@���˒�@����L	��tq����KG��|	7m�}�?�Uv�)�����+��r ��}�^��\�_J	C�ݽ�t�r9L]A�|�`o���`EC���%�Q߆LT�c���S�~�B!�L���{8Hk��m����ga:`�<�=��P��Ƭ82��gU*�_zo$4t�{˨���٦�����zŠ
������f�/�7\�&<A��e^ڜ �u�0�J
���GI.9��j����P��pHcw���D`Z7��4-(�^�0Ȟ_��6���$2�X3Ƿ��O�,_0?=���7�eՂ=}���y��ΥCa3���� �D2���*|K�6�<B��f����[!�ڋ���rgc<5)j8?{
���e:���9����S��L�w��o=&}�q	�S�h�|*�ۭ1�<�V��"�P��i������u7�9�
�yB�Y�J*���P�	�Ll����}�L'���+^~ ���3\�R����C�+�������K�4~d�+5��u��r'�#B�ީQX �j��'�Ex�)w%��
>F�>�Lc�%0���=�Y)h&w�uu=�{����ȩXaO<ad�3$�Y���Bp�Op}pY�E��7L�c���[΄{Q��|-YU�UD�6"=!I��>-��[;_��j��;���ySQ�����o��u�l��u="�6�"B�kkP�i�5�~��I�DI�U�`Ȗ�-u/)��R���#Wps錪�PuK3��y�\���:J�Om��.�
���_�|�St��d\'6D��KK��+���
?W��|+��vg|}����y+��
�(J�V}�ϯ��W�"m���s��w�e�'�C��>��,/�7ִ�hħT�|�H0c8$�� �6k�#^ay5��rc���'�d�Z���<�Ɲ+�U.B �T5�PXW��Eo�D�J$ "��o@���p�Rwi%��R������u�o����ų���{ƥ�捨�LP��Y��5[���䝐x��{�m>�?{��(gN}�:kt�-V�͗�I��#�l�P]���Љ�AE�B/墕I���ϳB�x'3�9e��]����]JBS��>#+��0{�	p���9�����U>�Q�+���
D%k�܈��#&׌�����o��9V����g0�?�jr���aA���2'����Ѓ�SP��7y�ݷ�Ɋ��o"�%!.���`k�!;wԂJ�Vj�+)vȲ5k���g�
�i_�/�??��쫐�Pϭ����b�=�qr��uʳ��4	tv����h���j�����;��.�_j�̓��tz�ze��Yk��s}vp(�����N�r��t����Œ%��6�"�e>$2]���J5�q�F��eU���H�:��.�n��~j2=�+X
H��8���W;�jh�Bf,�뛽��i�����Ni�1�9"�׭a>)�����DK�'�X*���j�^�	9D}�X��jy�&so�	SǾ|�Y�#8��[��-��������9l������ �X2:��U"צ����_g��u%����;^05�o�:���#y�e`����U��ƃ����J\ ������T\����UK���H�e����o���ͤ�nH���F��p����t�c�U�X�[��n)(�5��y�^�J�!��]�Z��|H��B
�B���^A�&>�5LM�B��/>Lw��fB��g�[^�.i��\����	/�%`��F���c=ڦށ��h��_�9����D�ƥ#lJ����=�*�QI\��Y��c�fʾ핪�����}��J���Gx�r��@�G��	Wh�"�fW����EC�������62�l�e����������˅ �������;q;'�u��� �ɷ?$U}�����,�c�Ȫ�6�P������H����A�Z��L�0D�ǘW�jc�5��}bq�;)����H������K�42d����0�y��!ݳ��=�G�y�,����WopjxFI�W~�P�u��>���ã�迭[,�ϑMW�@�I��r&���#{���iu�t��t���8��*�ef��r��Y��o$���~����C��ʶ�x&������7*y�D����MJ����M`�[_����,4��b	)9M�n�LW���s���O�h:��-Y�P�ifޛ��&��.-�^|�����:w%o1�~i�_��|�I�k��:H�/K��x�X�%�S���-[,�.�D�ͣ�8:&��g^�P"z���D�sь�'f�[GpA�������-~��ǀ�'��/`.�j�F�{L��Tz��6l�̊�?سy�}}���<��*�"���]�)Ly�
u����V6�g��W���r���Z�����M<�g�������q���G�\D�8	��0�C�HJ�@��PF�/��\�V�H�>���Z۞,弰~�f�rxfWL��O3*\(Nh��[����% � ^{�d9�@u��
�P�J�����$��ez�&çi�	�?�*�"mƅ��HՈsS����������+2_��N2�}#eB�".��Ӗ�gj{��oVP� s��{>�t����ۉKbb!8�+� W��T�����>ԖrOLյ������̴_�e����)�M�kL�����U�rÑB(S<�-� H���ߛ����"�ǈ��e��z�yVC��A0��+e<K������u��c"���wsw�
�0����]�̀a��M6G	+W}��h4O��-��ܠ0	���bÀ���,׭�;]q
R��� �^��k䷆�P4��"q<�H�V<�#���OT��N̠�n?Т0��I���p�͵��t�S>a�=I5=�4)=�E�KnlJ�b\@V���D�n��eW88�S!I-�s�,w1`N������~H�:\��ʅ�_o�q�MVN;��o�1%�t�4��~�7��7���8�e<�ݾvC�}e�IU.NVYz(d^�Swwt�Q�o�(Y��8�����������z#�΃�ZK�q�7�����8�����F�'����(�*4k�&|�f��.���0�������)O[(@�ӹ�����{!�I��@�!an��R��fc�YVg��pދ=j���᥋�G���Pp�`.J�=Tf���
��_�*������%V�MFx�lm��.T��@P@�Mb�������\�u\]��!�j?Ew2���_�F�����N�<��퀕H�w�sʂ��-[��%���&���l�0�
wG\8$ҏ>�U=c���>B�~��y�)�+$?�6^7��������'��>mV����aj��.����Ml�6_��(�F�V�ZS�+�U�ӌ�2�T���Vȋɀ�:T�etǜ*���;�܉��?�MF{����#�4ڿ葬�ڿ �_ G��}N����ۗw����_�#��]i�g	�dP<����3�C7���r���D����)��**i�1���;0�Ѵ��j���<�b%�n'��G&���]TD9�4&�ğ�ͩƷb�ݲ��6�,����V~�[����@�)U���1<�����	�����C���ήs�E���1�K�Г�����4�]HRڌ�^{k��i�V��4��7�'n��8�+b���^����	��S2;w��un�{[E$. S ��_�W���:�?�f�=�_���h�2Iv�.�/�9�Q�vt`&��`��!�f�C(�*1�eX�l3|��$�qͫ~�W��M���`u�(6K��A��xI���?��XT������[���"�,,�ؚ�/��*��I ���"��(w*��rbr���4}f`�3[:o&��gWJ*�UvCR@m�>^�䌫%3\g;��b����5���֢@���0u���R�|�{U2���#S��G�^Qdub�_@c�rW�A~�O���n%�{\Z���\FF7=n�	�Z�@חj��?)�}�	�fǞ)�~Cj�K��_U�K�<��V����|��f��1�\!_%_%���r�❅9F_���T"Ļ�&�:u�dd-8�!J��^���!Ğٺd���(�m���=%ӏ�u|¹ݥC,x�_~�83bH_�¥�	��&����$M�ai����o�Tg�Q��)��Mۢ��_�C_OC^�(��o8�Z0�4��Y(���j_�]'jX�F3�܊�m��	��T�=�'�	�4y*|"����T&T/|Y���K��oׯ�	���ȼ�Y�A-Y�U=D�v�<�z�����-Em���^nc_�| ���M�����}�8?�Y��8y�O���g��hú��B�X�*B��~@�+l��s��������l]U�fn| ��y<0�t��?�6K��d������v���Wb�Z��]WR��aV������A�h�*�/!sU��#�o���#�K*�ŗ�N�v�Val���5�L�)�dt�"i�~�]+�=����ۊa�S�me0J�\yg�j��2�+⛺���!*��~q��ж�u�v~��j�K���e"9�C��[�3��_@�?��?e���S��?.5ug�	�� q�H	9�%��o8ko�UcAµf��4g�EZ$�\�G�ҌO�gZ]۽�&Li�]���cRp��k*?у��:��z��Hc�l -�ܝz�ЯMN��&@D�Lc���t�.�q��Ǜ��@�G$O��/�A���P��3�d��$Iq���%ʠ�v�BzO
�n�i��p4�������iH^$��B͂�S�
W�Ⴞ���:���&�!���ZS;���Xh�I�Y�S��Ci�F�f�y��y�n⧖u����T:'0I�Q>sG�MA�*qf�L�8� ��$�!�K+�4�Z�I��T򻨅�/�?� b�-�u���e�U���e��8��p����yZb(ˡb��h#]�~yW���Z,�i l^��
�.��Нi���$Y".Az4��H��۝�6��2�iI>��ӟ]���"���}��<V�O^ʁ62?V�iFw�B�r��{3���[v�l{II�sq��-�B�f�k�
�b��O�B�Y5��n8���~W��0g�/���:[N�te-�/��w6ΔKxI� 8L�U��;@R	��w������
�Z��?�F��x�+%�C->:���aD���G��_���]�Kb��[��,�s��Q�FYv5��vK��Q�`��F�.�T�R�/;�%�%��� �Vx���$���Lc�)cV���lL��fНV7�Pq��O�;���Q��M���P$C��Vc�-�c8��x�n�� j�C�[~'�Y��В���C�pk~>�����v��V�~f��ըZ"��}�NyuX�n���+3>7D����D4!@�Y�1���7��Jȋ@d?�@hZ,�l���%~��M�� ��i{��'�G��uyDQ#���;J	l2�)� Ō�&�n����6��R3��+��w�m�~f#6k���S��E�F<d������� 3]~s#��NC���R��Q
�w��������*4WU�yi�p�R8�P���'i�;L���ۖ�E	y���8���	t����:�4�,+�7�!P&��) *���(�[o�`�M��flj�-������d_������оe��
�nsy�5��U��ޢ�#40X1j)~�E�]�4�N���t�|M�M񤵈0"�t�.�Liܟ�t�M�Q�G���6v܅��Ԩ�Vdh��%Υ�=w�~����U��9�n��r�����6�Cj�_����}���{(D>W�	|h\�т����l 8{���&���z|���1���A�r��p��O��̊����^'�E�����h���2r�Ռ���wr�lB���
|6��	e�� Ϫ�)���t�t�Ch��̝R�e��#"�y�;w�e
�b(������5H���1�r�wl`Ʊ%!C�Lԃ�c�^ �=��p�l���<s������G��2f%Q��ahWoN�@e܍�؁]ٗ���MB�����d���փ**m;n��V��� v�Y�T�����e��=H�]-��,2���7��ѝG�;���VG�7V�C�a��;��ޥ�eՉ1k�(�Τ��(v�W��Z��p�)N����P��J$Hc��Q�d.�H�6��D��9cN�>�8����aw��l���wmV�,�h7Ӽ�#L����n������ya쟼@��s����=���l�"lK])9k�}EN����"���g����e�q�P�����<+N�Z�ӧ7�	���.Mm�$.g'��$�`���za��������b���˦�ZK�X�ϩ�뷄޾��\-�����@������ׅ�ۇ�A�V��o�}�X)X�IkT��zg�h)��i��9�E$5�%�g璯�9�B�Cj�߾�������>p���e����_��k���*?q��g\ެ��+��i޳U�R8�����h��>L�O�~�{���g(T��q��B복���"P�*�%���WknhFǜ+sQ�8��v�Ja%t�1+���Xśo���6�j�y�H�ټ鹙�ـ�/� �h� ���;N/���Ղ����d1�땅�ӪȩO0H*T����o��M7i���i�/�{�&k)p��=� N��
�y���2+���~�Z��g������i�(�-ښ�n�������5ID�^�]`���S�$%���W��ȃ���ۡ�T�/��6.̺Q�"k��pR�_}����f|ߩ�n�(�'�Q�͚격�@�����,��R�O���$��k�fzK��`��bw��Q�%�y�I�������pR0���~��J]Ϊ:ܵ�&gj�jd�U���;��Tok��hދ�Ol�l��ڇ8��� X}q[�a��K�j�����E9	q��t>8��@�r�Jw�ګ� ��&�Y��R����!F���,����m��^ D*Z��(3d�윤��y'Q�<���v˥Y���Mq[�`7��Ks�v�2��1�I��3.�0ąh����;}�6�`�I���3ԝ�/�S�,���!mO�h��Q�O�E*��<M�QTu�$�(B�i��Oy�q�������]��OǄ�VT�msH�6 �h���@Z���0���#���ތ�'3�ʠ�l5��IR��������Y��������I�X"��آmw"|^�7���Z�]}L�|wC�9�M���»��|STn�cJ>`�\ɔfi��%Ӿ0]Q|p��quX;������,�����U�})Ia���km�/6���1��x��_�tW�-���,$l7F$�"�C�Nx���~G�=�APn��]�;Tߵ�TQ����"���~m'�o=����rV� .�o�Zd��Mo7�*��URi.��z��7k�a9�4���9P�ϣY�w����_7���QS�l.K���!�b:}��V�Ir�O��3a��e��M�Z���Z�ŭE�D&?�D-v��j��+P�19_6!�ɩ?Ҡ��!*'9�e�u�ӌ���&�����9�3�w�I�M�/;ux�R�>�c�Zn6xRwa�����!<��P�a����T��Z��Ql��Rʒ�ܦ��8��.ۮZk�o�	��>F�o�c�4b^$bq�/@�P%�'�������S��W!7_K�C5;lo\�7�i�����]Kr��A.6Q����Wj=w%����^u� ӻ�|{Πg���j8���k�w��
����{���K5�qp���l����w�V�XFS02�FO�!eS�:�_
JW��n�>r7���x��1��G[��y�'��/�B
����<��q�����:q�(j��c�	�mlD>$���h-�g�&�O+�2A��xY�)���}R�J�S��˛�ʋ��g���2%# Mi��ϔMi�R.vl�g�ȂF��؇���s���?@郅
`��T�t�3b?���^K��-Z��_h�L*M��P�a�� �(�t5�������ܡK���y����16k�#s�<vݕ=J..��#[�$)�.���,.{����_p%MP��5�^�U�\ݎ܏�����hש��W��f��y Ԓ�^C)��B�B��9�n����K��/�-���+�����m%�6#�� nt�Y���3N��.W�L�t]�JQ^�)�vq��Kj�-9�����v	�P��LL����m���L�ٕ3n喟�80�ܖe��"���a�@�䦘��-d��5o�?�d}aÐ�nrZ�K25LLL�I@5����ܟ���x���1{	�:��n#���w<���"뺳�g�ّ���l�sDve���;��e�MD���$EQ�R�ӷ(կߟ�����3ޯ���y��o)�=�V�'F�B�<�U�	3d]��}|4I�Éݗص�$w��|�����wҼ��
I��I�l�C�.O`r��n��Ѿr6~!\�r)��C�x�o$�Ý`���#�HE5'a ��tprf���.wbl(-+��z�0�/SpA����P��W�z��{�86<8w�4.�9�WwW�VG��]��jea��q1LM��x�����c�4���L޺{�AC���;����6[e�}�\��Q����#�1m
�%M��ћ����-ެa2򚍡������W�,a����A{�`�]Y�Q�3�ԍJ���Ƀg'P:꿛�뵦 ��+�|�j"֜5�bռ�b��t�G�{���߉�r��D�j�5�ǟ��PDq#@�[�D�ۙTs\��t�ɡ>I��C��*���,zQs���H��ʘ��|Ԣ:׳,�乪}e���_0Ev���ʐ^�Z~�+CE�4��gn(&esǅnΖ21��l��`����DW���W,y��u��Y�I���X��δ������N�_�ή��`z�a�"�cR�	�x�]C:t��m"��լ���`��q��rZ���F�	s�ėe���4TVr����a�#����n�ߠ����۰L�*��fO~3�y
Ѯ�
�Ӗ=�;RV�$L.yZ�����Rg��`��'c
�D�D�_*�e��jf =�+l�u(W�w�k�d�?��nzhg��'V5�s���L���_�4Nє�ˠ��v�8���ű��%�5�3�o���!�{>J�5)c�mǉ�lb�����<�S~Sޅ�R�u\���?0%���|~�ن�t}~�@�泒���nB�y�td`s/*Q��d�>uR�Bs�Tyj�:���r�:VW�2Sk�+��FТ����Rr�h'�!
�	�Uȹ����L����~hM��t^
��J�:̦���<pJ��"����s�Ţ�һ�N�`���GVᖾ�<m�a:�A�!s�c�#p'����ʐ��@&&�7�g��{r�2����2�>�!���:`���G�uE�M���;��p_�k��L-Q��9'�N�by/*\"Lܝ�ؘ"����@=c�� >ΰ �y�m����uG��>�¿����-7|WB��%�ǻ]����!|�Z����o$q��L����U;�ɸT�0��Zo�S�z� �)	�b,v�L9M��N�t����j{�Qg��4� /eG�s�CUl�,=E����(-���|�á��B�ne���>����EW[�����~Sk��PǨL5pd�Q�=:��QѶ�@�KGM��Wt�P��q��o���9og��j_�ȯ���U���iL�	����0>/Զ��z%s�<�[�?L����=z��  ��Z쿮>������
��"
��������D��q
gq�Ϸ�Wю�lE6q����z�Y��	qf�*�E'���M.%"��$����5U��-��Fާt鸎H��7ɇ�Y����:͊�<(6B�Y�2�xE���\;9^x>]�|j�[V�D���5JR5�I^u�=Q@C�ɭ��x��[�+�� ��.�p����|9�/A�8$j�/�)��te�T�
j�<�#0�	�����`�Y?�y����7�����
�� �+w��!���g�f���H�B�R2��*I�q���N�vL1���p���&���H4�q�jU�=GPV���e*���	����w��y�=�a��������ζ`{`"�츞�|!�}i�e�FtەȔ��p=�u:��IF������'�����2,�չD�YY�%	R_�y�
���3ު,�����ɉ��c5�׼�2�#�ɍ/II�����k�-u�⟄�]�O��zu֓�]�\��(��	�o;2K����eom��D�{���t���}K�
U� �^�c�%�
X�X	�_��r^�!����d}
$®�����^����X�*��:�Kc9�nV<��8�I��0�%u?5�8�ך齿�?��9�}�/� ����ϒ���ڬ=�@��՚�]����m*�;Sˮh�z6!EaE�ɑ�r�7��@җ8�(�g�ߟ�p�v^�Cw:�=�W��WsP�mϏ,lJU&�b�o�}�[g�m2�`x-4����<sA�e(����'}E�2&u	ZX��(&��+)Ɋ�:چp[`��35R�o�8�����4`��� �<�4{e����t���F�Ϊ�0a�?�?�ۜ`A�Y�ΰ����A:'?��������ws�c�;
�w2`3����l�����վ������߁����8���G����.%�����y���1�8�u�u�6%{K��9����LѸmI?���V�Z7���H6�R���s�����c�5�^ʠ��=歹��E++�y/J�k4β��EY�����N��7r�|=U�j���w&��J�{QqNY}���Le'j^��'C�Ǒ�bp�s_�]�fRH�2�!i�`Ko�>gr� hYT��P�z�f��5"���"���lq�����^�_�?Pu:'��������`�n���{��Sq�5A̺�C+�gc�g���8j>��8%+��Ѧ�'��X`�C���b�bܨ�4{�of����,���v�\Ł%����M?���߇'��:���^�d������	ߥ��2r���[~��;��ޫKTz�?j�YXM�}����%�źo��͡\�͡*h�K�<�/#�k���D��o;ϒʆ�\�0;>֫�K��!��Q."�*����'8���\���	V�ka�G{'#!<����ޅv��DSKĭ���^���� a�itw�G��&���	���Ě����}ƻx'��G�b��ގM҇�hM�a��ｎ)��M�0f;dAЌ-��9(��k#̜w�9O;����ｴ���a���~U�M�
S��l	m9$�Ga�x����w�������m�d%EK���h~AK�x�m�W��K���;��ഇ؇2�L[�4��l������f�B{�9s��?�?9��Y�: �ؓS'�i ��*S��g�H���'�O�c��4ǟ�Eo��e����){�wX�x�x��YyD߫&�+�5 �B����fu[�U���'7����o�=�Ut��W�(��:����AY�ғ��%�*�cv��td	�/�T/��eMݪ�t�y���(~���=ģ��+������!F�Y ��m�V�t���~��o7�b�|G���#�d����(�N9;�2KUs�2 ?����V�lZH:�������]3���jH΀B�mO���A�(����$rKٲg/_��|��@�� ���k�(\�i�AQ��y4��D�Ա��h:} w�պ�:�]�1m^&��H��r����A��!]
��VکfP�_�fǧ�/�j��qCR��m{����^�Z�����CeF�.��9���P�2�8�,
3�� �������e!�}�y���c�Y%�3��/�ܬ��`�3z��V;NI!��n;&�}���u�pv������a�c�}����eSx
��L�=���ZRz���MɬYc��FJiįh�m�/Xg�������r����^�J�����X��D��Z������j�mV-վ3�*Q ������Օ�����Ո	/�ޗo[aK�%��7Q��/���H�+���d��m ��l+(�Y	���A��vW��$�� ^��@�;m������z\����yQ셶����1�^��$��*�8u��L5��a��:&~��pL Z�N).�^:��}��v�֭`�#�a��Y� Zj��l6/��
�#v�G�X^s��fsG��<�Y����i���R]��~U���:�S� �q3�����BEo2�C-
�]�9ZE�e{�E�D���P��x��k_	�8Q��%�D��1�!���u:�H+���_�J�~�9�KƆ枆���tFQR��\���d�*E%*�я8��4�ln�4Ly�p�=�u����*%�'~y>]̡ ���.�xS����@vң�P����W��X�k.��A���n!MLC墉����X,�W��$D�V����^�a��נ1z���X,�J`���)�r�p�~��##�*���k����'��-���%�4|UjV��}Ω��`�S�+G�YI��#[��&��"W��j���O�)���3����W����8F0��~i� yK�	��F�.04%�5� �(k�W?�i�UX��hr<�C�v�ܜY�c��+o>��C�P���z�i�f2EɌ����L����d�k��7`�OD;_��=�X5n��J3����dx\Ax���5�K����ڣࣶ[�`?�k(ϼ��8������j�[�����o;^�Or$�	�׉Ai��Yh�l��kl%څ�7�ꐃ�g��21c*c�l�FioŢ� m�RÇ��b�J��{��[��?�Y�A�3*����8�$������f<3$�A�3X^��H�-'�v4G�6JiSS�[/+�1�%�#Z۾N��_Ap>Wo���\"�IZ��T�5TE�������V�4^:I)�y��B��6<�9j�Ԩʻ}i�����f\XY�|�no�p%=��Z����ŵ4$p58?ܝvA܁f1�������
�?_d�[�u��p!�b ?h�7��nT:����������!����� Ց���[�����5e����_��*�}�i�+�0���Qh�(dVzaXw I���J�7��[��e�J'�i���%Q�/S���X#����ŵ8�f�z�8l5�jkN���S�_ ����A����:^7����ġ�{y���7��a��L�޽v$��5�)>�<�`k�5���t/w!�Mt�P�I�,09F�ɰ��wyB����_�/6&��	DGQ4W3��t��d,߹>�\0�j��S(z�2n�Ú�(�|#�Ҧ���*�MV-u(H�WP��$���<�t�}2����A�jr��Z�}�e���'��,	�&l������<Q��p�N4�9�$[����%���cq*b]�[I�k�`	�d�ޗ?���r����7�x�-�
�Iw�ϔ���V8ʞW�<���?C����M���w�TD�o�A�;����f\�L���b��7�O7F�%�a��b�_Z\p������nȋ� ���3�b5Oh��	�Į�p���qB=���,]���/N��=��l(Sdk��u�pe&�"��+���{w|y,/�ЩQ�S�x�Ť&[�P�yh|�"���XqT�`�yr��'Rz��TT�q/��X_L�?�2�D�R�-�eU�q6�'<�F���"����s��	�Xx|��������y����4�S�; kH�pJ�kgkB����yX���Y1o7�9�JƱ����
[��;{����H��F���Ұ���κ _��,��A�'���L����oU�����q4��N	��ٳIm/.I۽p�E)�����l�K�c���R*n�^��;q��TR�Mַ_tt�"�]7�����`L����}��[�|��eH�m�H	��|��q<-���˞]��'Xu�UI`�d����e0������^\�r��K�%�����	L��y��5��3����oZ��n�~�M�g*ǻ���dB�|j@U%P�M-X�c���[Cj\��GUT�w�`�b�TϙL����P�	w��9Rԋ����0.���[ڨ�:S�>��l�����̐��e��K2�Ǻ_!+��7�	�9��̔�Z������v
��8j����^��:HW�Z@�2E'�¼I&A���(c2�(�z���x^Og�"�d5�)����&w�F��D�#��3X �څ�_�,r�\WA��e�g�\��&��eu@~Vm�ѡmZ�^�L��M=��ߢ� �֧�KYu�aM�e��Z��h�����E�o�K�ؕ$匧�T&=����Pb��܏M��MK��XdW�:m�r �(�/"_� 3֙2i���[�,%�!��P,�ң��K�[��#3��6aK������R`�����d>ca�$�u7A�3W�5ĩ�Ζi��R��t��0���\E��+RkE\�=n��Y��k	�3�g7J��(�7̌�%.���NX}_�\����{��1��� r�X� �D�_�oW�3~��<&� <�pz�﷗�N����vF�,R�D�X�

��Af��)���˴E]3�<a{������].n�۵E���N�J��Ũ����ݧ�?��CK������4�
����^"��!��cR�?J�G�5��C��]�[ˡ���1{ ̈�i�lӖh_�ȱk?kC�X�)y��c]��j�ߢt��8���ӊ��񨾻(L�m�B�-&�F8����3P�%��'�2QLb�pzL:+j�4��FZM�[�|.����?�rs4��(TC>�|0;|��q�ZF� ��K��. �J^g"`��V���(�Gy��A��(����٢bOO�ԡR6��{~,�8�?��:޵��0��68���2��5O���Y�hf��u�G��gv0�,��f^��X���D'1�W,�y��6@e~{}���|��y�˼�|�?����a�R[�[A�W��e�%���v��R��.��t�>����!^�Z���'��[�����)GӴ�+쇾��˱�2?�|U�؋֫��U��2�m�E�]�&��Y�mչ�u�(s{;1�!.l��f�=f�8��,^�n	�V{��f�=�Q�珪YD�t��{�[~?tV������F��' �e��P���[+��N���3@ݎ��ި�]����K���HP�����mg�	�JQ�{ I�L�W-*��	�p� /�#�<j�(3VVx�-�=�6&���rf����t�ʂ�n�LDr|>Թ�dK��i���͒�@+��zMh��:N�O�"?z�CY�<t��y��]���C-T�撺I�
�%f�t�!�8��k<M@�Z�W��ٍ�Z�{n�F� �[hG[�V�y����Q��s���M���ݳI��z{�pd�+�o�3�mV*soj�րo	ӭ���]����c����*���ظ�u�a�!~w��߭��V�eq���Kj�e���.שf��x��A�_ȝ�m@-v��a���<U�2��_'��>����J^�<^����^8S���Zdݫ���ֿ?gjS��#�gt�`����1���M+G"1+!�dB ����-�ܮ��
U�<��,�~���Mԃ�� �U#&���ܑ��כֿ���qPܷ�7O\��^�y�?�<��Bn�д���ktfK�1ұ��&���7��ҥ+����B�Mb�DYx�M0��QϬV�f�󡃐{�_���	��h[}�?��P���Ew�?3K�޺QS�Z��;ޓ'0Z��q�v]�X+?��ш�"H�3�]�ԃ��j�	R�^��wz�Ŷ�݋�u]�4��0ۑK����$I��Kf�g�?�M����OP��J�l�����']߃�����τ�n�������h�e�vz�Cs����+�E-�4J�ș:7Z���|���H�忠����>D�W O����©(TL�2�u��Ŭ����̭���@���EG���gu0���e?�!ɝgS�q�D�/��4׏+I�H�4��k;���;EN+���|�n�ah�=�<�H��S��H���(ᘓ��]�ζQ���Rd����H	"Y(�߄=�Oi��yM��eQ�c�'CO�;t��⏵"'%���=���U�r�B%Gi�M`�ϗ59�}����ї�=��e��$p`CGE�^�JpC�
���y������}B�ew�C�*�%�\�`���5�|z)Doּ5o��ڔ�&z׫��DN�#j�>icv���yΜCTv�4`�m�҂+×���m��a��Z~EF����_β��s/��q�ku��?���������'�ekRX3�m�k��I+�z�悿���Q��-͊�8ZJ�p�a}�ဟ�-�Lq/���W�u��[���á����o��ݛ��xp)S�Z�I(dV^��(��5�Vj�e	���-rb�!���pCDr˟#���k�<{"�lɦ<.��x~�yJ�EX��b��]��+fý�S�j,.�ԓ�l�2t������ޟD�TF%5���@Kxa'�����iyex���-�Qf�GءB7]�yrWZ曄R����{q��Qw��M��U�a�#f�-�U
d��&�ߌ��IQ� �A�xfF/t���q��0���y(oގXh�tuZ8��@Z5m���
m�Q�����e�xo����sC˦U�����Z��_�d�>������G�� Ǖ�I<���F�w�\��a���} ���D�tu����k�!V�����	7-�N�� �W��J�o�]<�b[ /c����@�Xe�"�ä� ������u�N�lu�#Ĺ#"&xoQZ~@�ջ�����lI���0[e� o�/��[�%F�?�:�V������\{�񸄽�T�׍��٤J�$'?cjY#�Snt�����G������[u�PT��8�ޟ�	oU���ujJ+��_'y�i���S�%q��$(���(,{H�BATz"�B��ִj��K���"�O��Pi�Q�8/O��V�SX��!+�f�-M0\�C��*�����b�)<(����0��bk�f�^Rh=�vOM���.��^d�ྰ�=��R����:�f�|�,P��}4;�c�[VZc"�i��xG?
��+ac�Ajb�<�)[ڷ�Q	ć<>$�e
yJ�i��i L.7�+�jcE��E�7"���-x��O�'r8Z����7��.��i��){ײ�᭔����u�Q2�Y�H��EłKqJl
5��Ą���l���)���~���<A�:1�h�cE�ѪYǷι��PNP>_ ϳ�^�
�p���^�"6	@�å�ݤ:�f^y��ei���G��F�F����@�>���"ܧ�Tms����QL�,���j��F����}z*�Bx���N'����3��>���A�}�בw쮺����{�NA��̟���7lP7���.�����	�l{�x
��h�e���Z1�T(��@K9�h��:mW�0���I�sB+,�p9��9ڷu��Ul5�J�,�΀�9Z� /�yR���ntw�	�`�9z��⑄�<����۬O��fv=׉!W����T�p�b?�p{P�<%gy����6qƒd��q#����qRl\�L���}��)��P�f�30�`f��:�V��6�lG�2m4�73���p{����MHl;��'������f���cG���"l8¨�bK�`V����@��(-���@�߷��=r���MR��|�f��X�O���Z��BT���Y5.��/�
���(z
vT�5U�?\x�^�h��A�����d�@
�A<��ǟ�N���8�±~�!*�
D�3��w�TS�r�
٥�L��w�;�m����So}nl�f4�i3m����&�4�b~⑼n]G����'���a�Ny�]hcM��\ >�ٚ�J�ʤz��5V����O��.�9@e�1�"��+WW���5�@O�1Cf����4rl~�S�`���Cط��5Ń�1� OF]��Pگ���V!fOK����\��Eb�qJ�R�Y[�_ �pj�k�-!�e��60��D���5+�-�������7c/4����kԵ��y�P����$!���+O���&�<t1�����:\_���غL,�-�c���N��I��^��*5IK#J?mo9`�:~�������W��a�å�]�����_&MW��������w�����%�9F⎌c������J�_ѷ��S�n�Y�]eu��˥��H��V��$@�Arv������n�@l�����gĵr��bKE�Ѷz�Ew̹H�+|��r�.�I����(h��_�]��FÃ�ހw��"��'�ZO�Uv*���'b�7t7���1A�<��4���Y�4�ݳ�s#{p����X��[f�ǅ�ڷxw��S.��6d���w�q4����`���*�١�$��N����|(>��?���^ѥ�������G��^u�P�̷�9�F���̤���ܕ�81v�k��E�܅KDbkiH�6��Q��T��n��؜�81�X0[d+�����D����&,R�P(q=���[̾�X0������=~�1SS8E��5�g�muze�� ��'�
���|[��[x���3p�^p�a��^JaI���e��0G�
s���C� ��Ͽx�]�~7�$
�#9�IծR��"��ʎ��^*��k>���Q��޽-f��� A���L��c�^G��W����{�	�oC��K�-��OM3�7�D��������p��}�K.�k���w�s���k:��L9|��q��A����1Z�dW�Ym�(�-�>�zO�D�V}�|��о�c	-?��� �@�6��U�ih�a\��{R��h�k�EH�e�d��� ��L^_��O$�ֳ��w���y~�.X��j�Ѡܟ󊿘vR����Z�ʗ߈����v�&�NJ��9�B�����A�U��H��C'٩�/Z�ti�:f��:���V5$���S(*�mf\��FW!;ú�Q����r_ʷX�oi8�7G�ZP�0
��K�P0p���~��m�&-М����^�!C7�'TK8O>nTQR�c���p�X�3��x�C���(V�=�g�6��Ҙ�V22e�˙\qd���iĀ��Y�FϿ��O��O���u���wYA�NB&�~H�S���DC��)ۆ�{�N"���>q�ܪu��L9��䓁�����l��?�7]S�T�1\*���3�nqc���U��-�"�N�h��;({/�6�HX߭������3��.�H�����¡Cf�@_?����E�!�-�ѯ
0p1l�Ä����Y=3:�w����з��Z��!�U��x��V�yo�*{�i}��,���G��ƛ��A��+���,y�}�z�\(.t�%4� ����#Om��n��Ƙ��܀�$v���;8����_r��u��`[�U�j�2��a`
�X�l��#�,�Ԭ�i��yl|���#.��ǮT���2��l��d~kVsp9+�eha7nD� 9=C���Vm�/�t@�n���X����]'��`�0n^�cm��|_줬�W`��ݙ�o�3W��b3�,����eW��G�@0�	�*�����|�����˳� �U��y }Ժ�^��J���;`7%��<��&�~s�����U�ǤSsr9�|�!��Oc�w,oJ�T��?ߵ�j_I��䷐\8=�֬�U+¶���X��Z��\�ً#���l��\\�з�U
'�FY$���2�����ʌ�NL��w=�������b~�{��]m� ���44�q�&�������n��FX̯��_j���DΡ����L�`h=�����f�+u� ?�ۀ��*"~�8k�y*<���͋L�Yz�s����n.�F�#��0w��s�3��3��%�가E�`��O�^^+p�pV"�D%#��TL��.p��X�� xw._��d���i>Ӆ��wlC���� }��2�����P �φ��;���V�(�O.\���@���^~ !������h)�11�P+w�=*�'8���Ɵ"(�ula;:�F�z����1\!7���{�z���r!)�����Qʬ�
-,_��m�����c�q^� r
(Fa",<��kE���[d�Z�׈��kƹ��0�ɷ��p�;Y ����i��N� ���X�)�փ>���<��V�o
� ~��cy�1x�M;?����w�/�n233}�	s������1��	ӗ�,�����g���BX�*U�<@=�ƺ"�Ԝ1]d�r�U��ϰN��_q7�ڊ�Z?g���4T�mk �a�$0�J�r��o�,EIg��N�����UH^��&��,�ICZ�.������W��#�|,��u�^'���c�.\FW3�gK��$���;tӷ�s�u}p!��;�c�]g�� �S+����ס�-깛V�C%(�U�"�`��9�[?��]m%��^G#GJ,	��VG�|�Y��a��=�L�{���7���4�0kHe�t{zdo]N�u��x�s��rZ�D��6Pr��Q�|�5����mlc�*[�@�Q�v����O���"u߈+۱�Y�N�H	��s/�N�)ڝ/B/�+���w�����q� l39N �X��5�ڻ5�����|&"�x|�*�{&W^ɋ�[���p��q�Fc�����y��	�^���<�)�������>3uϵ۱�ž�\�Ⱦ�pė75c�kV,��-�fʡ��}�_Ӟ�]�3e�r��_G�{�>TΞ����C�^>s�B�U�P38�����J�c�P"��֝�����C�$�{��F�Pղx���(*��vª>�����c(�gd��J�)�*�سCT�/qwϲ�W�n�k�"ה'�E='4����E:z�m��wu��n��KP,��e;8*����@�/�e�&�h}~O� �dN��E��+�a�Ê���>�^�����0q�L�:F
��Tn^)��b��z1 .l�����u�h;}�+@#&����膗��Ir�.�q�> |�B�/A��]c�X`¼P����G�����F�ѕ�p���\]v{ ̧U���P4��R�ϒ��t��y�OW��ܱB�m��*��ֶtj�﹌z|�y�S؝i��k����+�h�%.�]�;����;)���޶���W�8��˄��=��,+w��>X��֥,�5��,z$e��S0x���ҝ�)�ڽ�I�
[�-dg��B�"r�tn�X���F�q��Ɏ�����m,��d��%��-x�bJ�&(��-�����e�bn�D?-���\�B�G����
�o��_�kr�J5H�աB��d�����5M��7z�W���X]�5��Q��N�,Po���wk;x��g��|u��~�'͏�x��F�������2(CT�ז_�V�����]���.�ٜ�=�"]���:��cIy�԰��~QB�/A}eU/��H�]zMM��>0��Ξ^3�$luy����z��$��g�7�c<�=Ѫ����
 ����y҉ǣ�*��&��u#���57:>��Z�HN�Wj�
�S��tLͺ���_���m�oM���SV�[���m����La�\LE��۶,��P����G2��Co�&��� ���>_M��ъL�Њ���D�]No����%t@����q����@����YS�(���F��.}�������� ��i���"=��_�D��2g���\-��6�g�n�.F?Jh_1.����s���.��Qo�q��eR�X	���4�&��)���B���igP��oq����1�;����(<D�~/E�l�����ҥp��r~�m�b�LHC� �D^�Y��Yt��3-D�a��� hw���n��{�a>��<���<�?;�є�0-I/��/���k;[yŋI��\�4��s���@��R�>3�Ņ�b���i��X�Ô[�ҍNc��m�}d�\������w��~ G@�Ă�� Bq$����#���Ey�xQ��%AZ3Fx_�k��M�+��?�/��z����P�}�X��#E�+-���y�x6�\%��fٶHg��hd6m>�9{�4����q�z����)\/C��:�a���L�A~�)X��D�DY�k��nC�����3��&�!3��|oF��D��3�,�w��J�-CU���>��+(���sb����L!�r.���c`nn�����% ��Q�A��2�rZ�:^6q��4SU?H���Փ1ox��pu���#�γ����"�Uϼ�-
�$n�`�;�>�K߮���3���T�C���Ky���/�7N���o+��ܴc����~������K��$1��(��@�xh�̮���Ap��ݳ?�������;X��c?ἳ8=�p4�>.� ��H�����e��ͰF������NJ��J����ǥb��B��!zt����3y�����Z��D&�=�H��(��U�����9ʍf��^m�!s��sB��d$�'p��F԰�F�ΰ�H��WTN�C�~�"�8D��lrW������r���0�=y��g���"a3�0j�~�q��d嫇�ӏ��>�,+K����'
%���(�8ŇY:����I�ND&�J)��e,uYl:y.y���/G�^�?{����Y5��r��Q�F}������b�������q��?��S��dG��>�}R�*�J'5��z�ru'W�m/�Rw�P��/b�x�)l/|�3�K��z�=�	�V��,���R�r��Z{�>�5gɚ��MR��:a�/��T�_&��6 dFc~�����]o��UY��ΑB1��[�J4U�t�rN����s��27��֟^rY��()���YA����t�5�r���)b܍���'�r��M	<��(�[���)+��84�֒^����!� b�f�����&g=������\�<�&��r��kjzG����MK6�t��Ӛ)R$)��!��r�'w��V��i�??|����{ݼ���`����F�*�����\1�p#<�(G�#�y�m�)��&=E�'AaܓO�/LUp!�@�]s{�/�Cjg��mn!� hL9U~y�n�)i�w������E۞�t��ͪ���д|����O�I��3�����62D<���d�qS����WW�����v�O�J���̈8�)b�9���Mx��������Fb�T#�h���-@U`�}�V����~rV�4H�®���J����e�I?%�Gޅ;�q�x�a��|�ImEXgg�GG�;�-�`C�tHޯ��T��O�a(�'qk�N��-X0Ra˷V�S�����fǀ���zn���گ�W�f���m�f�4e�K!���7,x8��T�������ʨ�`Ii�֞�|ERQ5����U���}����O9�ۛ	Ũ��	K�ml@$�^[�v��i&>�:e	8J}���/p�'�h�=��&����"�·��vR�8�k��Y�NWs��� ஹÍӬ�Z�t�MbH6������ �Oz��Z���f� ��vgO�(�{�u�cŜ�$b�czA�C��>F7���V�It��h������я����1�����'O�"�)��-�2I�*v�>MLFBƬ��$_/kMQI#���wG�@���%�d7���S����=���`��M�f$��	���m�3|.����M��pITڲ��Ǥ��L��A�JMh�<X�\�r�5������}m�Ad��I�G��#���a��8t-�V�h�9΁ɦXY��CCI�ۭ`���f,�Վ
E>�����yt�^Z�>}Ԩ����{���ث�������.{�y���X'Rf��7�-���m��2��9�G��.�]���`�:�7U��c��v3H�� ="����c��$�i��2���H�K����oֽ&f��q�j�a��ul|
�� ��мP��a{��s�V�F@�R�u�E��������b`�G�̢�a�j����*D��$)��)qo�~�7VD�,��1'	ة����١�An��i�-��2p05��gAF�'9�lgt�M�u#�� Q1�'b8)�4CG|��F.=�7�4!���"�(������P�عf�F3��=
��j�a��?�gy�d!շp��8e����3��͡���o+V@1?$ο�eR	M�p�=�cooGkN;�%b^_��	?Mn��љf��T��%*۪�6(���[Z������ڿ0H? ن�T<#v����3W<Z�s��8��%�y�=jnǢ�ǻ=`r�B$n�F#+�����Fs�O'�Y�/��]L����o�myQO8��x�L�%�mXnf�&p�<�.�Fz���e�(�o�sN��~R
�8��2W��˶��@rx��w��d3a#��U��?R;�
�u�V�U�Y!w�t��/|#]�k	9�V������s�g�}�����S��qNs؜Y�gs63rH���$!�9l̙�sf�!"��9TE�bC�M��T߾��u?��z�����f�o}v�,(��O�AU�p���w�r&�x	a����Y��r��1̟�I�����\�8�q�D�,3��u/�J�tA��
�:	�� ��\-y&V7 yu��[�w�ݩ
���f�z��Ќ7��� �L=�[����d`;�ӶQb��$��$�\Vž�M����S���i�I�9�l(Zl��F�G�^���]r�j��P@����+�J���ӌ�]JΟ�Bg� �a�]�rE{���e"#!U:��,���Z�q��*���=|Yv�y���������.|&MfJJ��pb�D�+}��l��pV43��gw=����rm������h�#�t����9�Q���,��ɴs�}?!���(�>��ܸ�kv�L	@�y�{t��~U�ۊ\]��3P�BF�s�/�ټ_n!�n�`�KmNb�Gs�;���Yg_�n���b�M;C������4��-����g~t�/^�6|��wX�`�]����Z�ѣM�eYM�V⋔'7�k�����'�	}i�����.wC^�uٕ"Qy��τ�Oŏ�A-�������	~!�.`އ�'���k:�W�*�O}#����/�V�h�{v|��5q
��j�{��xV�3���^��+�^���at���3 ۪ ��v5L�:�v�#\ϣ��k+�3�M�ԧ?�g�?p�������LE��)$P�{0p"��>����Ϻ_��˩�?;�t\x��f3W���/^�B�m�nh�_��BJ[ډ�.�����U�?h�\$f���ޑ:�fC,�4�\ŝ/7*�������rj���8�ٹ�{�;/�S��_L�\͍�Ymv{Q7��K*�{E���z�����z^~'��@r4�,'�/�U:�+�P�t�I\�J�ż���>���}*�Pv��̆��H"^In5�s�����߮��O��~dR�i�l����|��F�m��κ��w��(��H;���b���_��tD]3KY��c	���Faɳ�ۢ׮l��QqɝuU�L�¤����W�{��e�a�_�S��oM�N�&;%@���۾*���ҍbw�o��"B�i�ْ�>��E\a��y�R�l��}���
�����������B(ڶ��'�U����Mu�ɇ����T"rx�Wf�Xp�	$oW^V&w&�� �$_U�P�S�O��h���-0�z[�Q"����Լv2،�K�l=`J6�Vu��Nũ�֛�̒1��q��&�Q�bjc���'�b�
�;l�Z�P���Ϣ��T�ð�n:�/[Ŀ���=����1NO�.D�\��ϫ0uT��)�y_o��%_n���1b�k�"q�a���Kg1���� ���vz�*Ӷ�Ӏ(Gt��T�IH���cO�*|�?-����6���w�	O6�4[ɟH��N�fi�L r�=�J�(%�a�IW*!8��U�C�Pj��p.S�˷���y	�4/_��A�����@�P�/a;���N�V�6־�4W���9���u	���֛��.R�/�hr�G�<��F�̾��)�fng�L�vw��I�N�f�ҝ�ʶ4ݾ]WsW�6�u{�na��, ��j�m1P��J�<��/4`���K]��"/~\���|#�~ז�6�{4:�а;�tRr.�g:��N�x��{�(�����e>��U�<}����1oj�m�_6�{�b�ݏ�%����Y�J��+*ٶFr1nG�i��p�&T��.���*rzֈ��_�*�x��!�H�f{U��3yb�f�����A��n�����"��gbV��������$�����:D0K���"����S���.<졵{��M���],X%���r���y~"i�&&�d�����A�֑:,�z)c�Y�ҿ	RN{z"��ߝ��ܖ~�),PK�6,�L}U���-¨�I��cx�u���L�����S>���~U���s���>Y�A^|C�g6&�W����<��aGe�Cq�|���E�����7 �G]m��j������N��������k���y����WU2�_C�1M�:��o��k�ZȬɾ�Ǔ�!�W�Ӻ-�*lϖ�Ɔ�T����K�8܎9F^� >�U{t��+�Ϟ��y����lĆN�
�[�cUg*�t.�Ʃ9e���G �h��n��{�	4|~*�O%����*8z�����4�|��:L]RoP>���ޥհ��G_��S\.i�,j�Sm��j�&u;y%�x�딣�O�w���J����]�ܼb����ϒd�-,޽֎J�+�7T��
��W�W��EI�ā�LB�iZ�,��&8�QP]Ö.��Qh�ك��!�`����ăC�L���"��s�<[����=RMuK��I����c��s,"��(Ux1�XZZPR
�)�P���\j4���~{�R�ý�7⼜(��t�*~&ʹnt1#����\f.��M�Wv��i+�1^�(�0��sWU�i�M�4�"!�rA!_���9i��鼫��U<�h�9oAϙ~����,s��<�x
�8@9-�����H�Nd4<��+1�Gi�f������x��ɟ"�ߏ�����m\�hA2���������˦/��"W(�y��g��jw`g�wL��T�,����Q�6��=�EK |NB�~���7��
_�(~�a���?of[7�u*���(�U���_{"�u�Bs�X_�8;���
���F��cKϑR�N�����X^J�(W\ό���66����O��n��{��;��.k�Ţ�W�>���T��kɉ� Z�����Ħ�����t[`�s2�90%`���&������|Ι�����rF��{Y����Ds������d��e1�����e�L������W3�y-�ޜ��`�Ond�s��'b�A���C)4ͣי��3���J�2�M��:_���ȑ����X$ �]k��[~Eq֍�9�La*q��<�,��b}��͓���R�!>�*���x?��d�_�,���D�@>IIe�4D=�X�K3�.4^j�d�5uY�{XjIc���ػ�o���.�¥Km�q'*<^t�1s*O*=��m{hh��;Z�;��PI���|��v�Ħ�}��@مG�0g��7EW-�Ա�#��U@����.❈վ6��Dw+6�#3<,�`����y�Ï�Kȝ����w������6�>��u�uc�<�SD:�а�O���=��1����G��c�D\3�����QŠ�}�Tm��͊�՟�%�V:�d�����ރ�dKeuר�:��ru�8]��HE�Q���S2Z+�g�
���3����)��a����z�˰2Dò��⫋7���.��N"kDU1E��x��;՚�K�RTQ������Qw��<v�3���2�]{�!ho�(`�I�v�b���&?nl[z�%Y��x��A
����D����)���d�߬��N�A��֘��ʮ>9�.��^+�Ug]�|��7�� l��O��}3e��)��Ai�aت�F�Ro΍J!<�)�<��K^/@904���}�O����q)���㿽^�u������%;/���^�T�b��w�X�3�X�ݖ�f!���C%y�G�L����lFd�rG�3���3�ku��P?�q����od��m�C��d�-�geo��ea�e5�G���ƞ� ��̓3|������-�P}rR��ޖXL�%��Zʄ�=Ҵ,��'m/��?�mU,I��!?��wG�T�^;w���ҡi�HE�H1���Ԯ3��q�DE�-L��eQLuɋM-��?���=�oA�[X_H��%�� ��#�f��w~̀�u�WK����Oż�H���g�@�cԘ�2�s�=�r�%� l��>W�MwA~}�">�j��梢~\� )�2�s;�.�ی5�;K,,x`�:�޴F�d4��$>�XV�ʖ5KQ�͵z��������D�{���.�|Ps����9�]�b8+�9��=������%HJ�s_�\��_�ְ��fZ��k������Mh���S�.e�"��-#�Ũ�"��0W���g��J���K��J��z#NK��~ҷ� �qb�
#�b5:s^v���g)��B���E�'�K羐t�xhc%��N�6m��Ԫ^��ul�,�^Fr�TQ���H}��;�[a~�"]�v�⎅��"U��U���fx�
ޗ5a�M�-��`��KC�)���n��@/H
ڳ�DL�쇰6`���@�[�qe�"�r����~��od��Ѫ"�yJ�2k���+H������%u�s�U�D�/S�;5WPb�}�j�(��?�V��O�~�Sw�T�e���c�'���iu,�ӭa������+)]�r�W"f���(?%z��xD�M���
���_>�}���Wό�����!^RQWZhY��Qˀ���t�Q,&��JPw���b��9z\^��g=r�+�v��4I�,P��E�n��8*5��T��}��!��.H����<�(��<�ޱ���e4Ò�Oa$o @�9�m+�~�R��� xi$Z��D�%�zؾ";Ye�F��b�%W�
i~$/�v/-"3�R����~����̟���~���%�Ě+w�Wu=��2"�<���_�Y��a�{�`�n����3�yB:w�z�wby~��`��a�c��ݑ�����+I�gBN/�p��7�tnB���l����o��%�l���|�}�vP��.:�ը9��V{.Y3��tK�$;����3��l1<W2�pt��ZT]���e�f�:�/�db�{><�@�!v�84�À��b	����a8;IB����������k탄C�4ؚr4=���2Z��R�aMM���A��:X�8�Oy�lk����i[���d�	t�5��l<' )�O���9� Uˮ7���u��ܔx���}<���uF�(�P9]���GR����m�����5-S�kw��ѐWQ��D�aLh�?m��>M�����R'M��l��I�ǀghx
�+�y�Ij}�=������Q�qSQ���*Ma�<!-D�(n*�O�4O͙����od�t����ߧ�h�)㞡%=�ޟ�'�M�����%��Wu��ә��������{�4B����Ys��I7K]N9\�
�qu��Y��BA�K�
8�����N!��y��Z9�86�
���e��H^b�aU P�nR���}$�|���O���Q"�!kE�I1�E�5��rϕ��
��0��>�G��Ѩ�ORL��[=_ԻT�G�[���nƌm��*��*�d83�������7��� �5d��:0�e����. ^Y�N�]*��~�蒙O׷�"�-rW���X���T~+q�6"��(R����'*0�tL��:�|���*��ag7H~J��}�k�81nDj�r,^u�&!��v=k M��"��f��,�E ��^�Wm�ő�t���xoB�"���_=�o�L��}��J[95���?V�z��·���հ�^+��Ӆ�_�/M�u�}��>O�|gSu��˜L�(�þ�V�
FN>�﯀�6/�H���>[��-ϫD�^
���G�]_��A�+`
P�2h����BG�+�H8)F���w#�51l|��������K��M�3�i�zNԞ���q#�ex#�«������-Ӵ"c«�d��g�ZІ����ȗ~$�U��D�ȡ�=��
Zߜ�v�ʒ��l"�����a�-�������hP��a��CL����A�p��6�'��������ԇ^/���bג~��Ƙ�s�0��8�w�sZ&�3���N�Թ�¼�be���^H����-��՟�:'lZ��T�H}��t�6z�� ���u�C�;ޭŔP��.�pE[�x^�]d���$���%�eX�T� �'��`ekd�~"��ס�y��QD�j��l��J���W���OP
OY�ۜ���P�����s��\�����KJ[�12��Y��ޮ�۰ݢ��������xD#�)f�ny4x������e��R��d��]U���C�Q��'�D^j����VZ|�v�Ռ"��(,���?q����yn^d�#��c������0E�mW�I�.�¢�����*��fϾ���d]��Ճ��)!�RH�aBsq���n���5P�Ko���dj¯�V��SAr���Q�k㗴�	��DQ�)x���d��䃹a�-Fʱ��5%m{�po0 J+p|��
1�(��ѐʅ��##��2+uR�+�:�����V�w<��[Ш�R)�7�+G�q��$+������h�u��B����F��h���D��yc'�8BI��Q���C��,BB)&~]Ui��q8P����n�џ(~� �e����aõ? �o=�ny�>ʱ�٘���Aa{ز�$cQ�0����`?���T�O�|x|��O1�.H�	��M���go���;��M��[�|pO6���:1� ~�H��N������*9=��:C��g c�s�m)���Rz�g�b�g��K&������ݫl���h��d]'���'�4��O�ۛ#^]ی�)�}��a�z_J�a��ߠې�K�3�����]�^kV(���)���t)��H��CO�K(9��@#��I�EI����m�}�x�z/M���?�Y煝��3���}����F-�b°-��������u�!WJ���1|Y�ru�sH���E�@���B��z�Je�'Bs\�1D"�������R��*��������P�'M���J��	O��(�
�|�ιç�f�=�]��5T�hϯZ��<7ߏ�����D�>B� E�+8W"N��R�<���$s����,��%����n��nr�9ć/���PVڸ]Ha�D���9��b�ʳ�8��������	�'���4u/�%��3*)s�׾;ӡ�KZ	�+�[�>$Տ�W>������P�lmL�����[Ȋl��hi����z!y�:�䗄��[���%_��H��!�̞ǝ������3�TN��V� 2�UE.�L�S����p�3o4�Kh���V���	�{�'�^>�k�;{����{R3�f�^ �2�u�k�ȷ�>�L�P���'WI�71�+;���W�a#/�=�e@�����Zi�k;j|��Мp-i���e��6�H����z��	j9El�*�zY=��?�Q��GSx��<���IM^(M��$G$�jرGL���@�j5m%�;\
�����x&&������3=�@��/���f	�����W���}#��M�ôE�j���L�k69��j������s�Uť�*��:��N�ӤɯQvM���]�H^� q�4W�h�J����_a#5������h���')^�05%�'L���(�,�9�1�|=�^U�?��Ih��ٻ�U'ϳ�9������R?�j:zQ�ĳ|O\1Я�w.���4Z�r�0㿾,]��3�|�D;��텆��&�wDQv���ȼR� O���G����������fi�/@����F�;�|��W��_�&����d��>0��:Ps;���~~~ز�&*R#�di���i�TEi$w��Uŋ2������:d��hUs�|�vL�Գ ���,X!��<���U�QP|��0I4��m��C�Z(����̢Ř�VĈ�A��!�?k��у����/K��9��"�"� �?(�i��k�`*��J|�,I9�-OTBJ�;�ɜ���2@m�MVa{��|�n��mP��Η�:-!2�<��UXp(�Τ�;��0�d:���Kg[��d�=|؅.U��Kй[TNك��#��<QgU��ms��#�6]����3Р�9\�:���h��Y=�Îl[� ����BL���|�A�=(�qUlW�K�Q�:'8�2�!b�ԣ��*��O)�jJ���+\���9U���>j����!L�̬|k7?:
��)C�jU��_�+ON��maAffɬ�s�	��=�������=G��_�1g�.�D	YT�D抣v��	Q��c��zwg|�Ӌ�Vɥ����M��rH$�"�㠱��Eꆈ���G��k�6���~!���Rx�!c�U��,xa�)>��c�x_��X��H��QkH�́n]Zy��cR �R��݄���S�T�QH��|4y�.��,�ͣJ��)5й[!!���"�M|*���3���Ӟ%*��W��U�9O|�W9:l��ߵ���4����W���s��w:rW��}����]D�6�j������c	��:�/�jS�3N*��6usA�B����E�T��?5�5Jf�I�Q�&����:������Rgś��B��В��e]~�N�bj̠��������)�3+@��2;���X���5#Iw؁٥��нpe���7�yZ��0qOI1�3����,�;�q���n\�/#�ڢ􇪣����Hd�rk��C(JC���~F��/پC���7R���-z�����a���XeRӚW�n���JY�wg�T��c��)'{^�ȖQB ��6o;�tk�f�`xX��}�8�ɡzOMm{�>d��"�����[�`�Ŗ�A��h���4�B]۸��"(�y�i���,Vx�K�Mͺ�����N�R��)c�kv���N��&Eڣee�g� ��RZ���!��'�+1���>��xok���s����J�`"3���\wR:#��ǅ��M��Eu�|(x�w_��3yL��ܯ`�_�"X2�_ӆ�/��o�\�yxG�̷�y�=�ѥ:�#I�Sk�����odp��
��eW|�#��H��~,���w��0�{�$'�֦�m���Ɛr��(���Vu96��N���S���C���b���[���dH�A��޵n�Td~�]�W���#���ly�ݞb"D��VF��U<+V�w�t��#y�T���&��J{(+{�"�G,?�U]Թ�Y��Î�C�c�$��	���A:t�Y�aY��(Ju���I9sp�S��I��ܢu�pā��.�W�v�ԋ�~�z|��1��G������l��S��{�Ŷ��eL�v���{)���ХCط ́zyqQ���*�@
��XE�5c��]G�iUΟ�ߴ��g,!,s�bh��]a'hi_��n�r��;O�����ڒ|Z���瀫ٔS�&��K���IE)�
_=��a��~��*HF9u��8��rVV��NO.�k�B�u�B���v=s7tI��/!��H"����\�霿l�r�NNO;]"TQ
?��>h�
s�'��Y�3��l���Q�C���P>�GaR綂W�yJ���m����#�]�
������k����kS�*N�[)t��Mx��}��a�X��?�I0�Q\&�q��v����%��ݷ��F%q��Y	"��*��h9���G-K��4�֪�#�:�~�W �>��gw��f��b�T���W��w����pM�+�"�g�ZFw���E\XD���E�q7��˻��g>��m4� |�z(����B"�{u��a�0���5Z��I���!C��c�D2��+��Kϙ�K��[�1)Of��s�CaL��ϷC����6�r$
5���6�~�?-��!ƉEӞ��k��t=�\c����ӓ�lp���6������i�������1��8�4`L5b9o&Q�y��D��ݑ���y4�KwUV1��V!�d���������l��-��{#,���#���,K�r�c-�Ɇ�ebԱ� �,��l�Dk)f����@��8H�	�J��\ �i�L����H�'כ8���� �烬g���H�џ�H,fiй�I�����晄8�{E��{|̑4�*��L�ý2�W���b�ةq��1���������|�k�i��c�ÞO�ñ��z^XW�n�2� b����j�<��*`�yWv;�Wsz͎�q�L�[���D��0�lK�*aw6O-$�iw�p����;�)��՝�h}P�l=�3��LW���Q.#�P��<���T�sT9��]��z(B����1�{pW�E�rWCkʵ����p�d8���F�Ң7/ۖA�g�
J���|�x�<�u����l
�>��we抙n2�wT��;%�)��8�h(!�����>CіӸF%�^��t�S�&5�o�(o_C]x��p��ٰ?u:�an%��m^��vN+�H!�uyEfj�Ȯ����<&k�A[m(7<�yw�w��ik*,�֦��}V�sO�h�
�����~�$�Q��"��H鿼��,Vu;��~D���||���Yȋx����E���<�=�ͦ����	��\
�xĹ%�$��i-�uj�I��d�YԶ�r��+@9J���g�nWY�>/Q9�w���  �����&Q��Svl{�i1?(&�����@�<��(�+9���;+2��v�w>�Y�/��k˅׵OB�m%��IX���^Z�Q��*�z���O��vƝ��t��Q���;X���cf;�����%���Tͥ�]����f��@�����E/���(��W�]�<3�V��R�������s|� �gGn.I�:iQ���ݰ�u�D��gU����zsD�M�5Ѕ_v�h>n�>Ԕ�(ﲿ�>��t?>GѬ$'+� .l�� f�IRaO��ڕm�� ����<o�q^��w�K]v(V��M�'��u8m7��́�2��+��$ľ%��ru,]E@��lb�[s�ZB9�ɦQ�nV9W��n��ɥ!��s[����VA�/9�_a����Tf��\Z�{��k���/g���o���y�X���F�޻-I0��V�Q���;��,��6n_W�by�)�ލ������b����AǍr\TOhP���FÝ��MN�I�@jSf���-�b^�T�ڐ=;�����&��1 1΀��ͭ�Gsa�9Rt�KC�",������%d{f˽6�}ީ�F��mv���L�=��0��2Y��w#�A��o^\�����$�9?^Oi��N9l�����U���2m*���
��˘A�$�s���9�Uh���/�.�7�m�0�Qheg�Ɣ9�ELgq�T�I��5�B ��˘ڲ�YH���	W��K}L#D���m;��;<��ϖ��d���2���Sh_��q��A�8a��eqQ�=��埴Y��J<������`i�q�/����]U���a��g�^o4P�(�L[���@���\���]xqޝpWyt���@�&��ji� �-�iUY�ҹj�Y|��#�WM�:��L������ecH&������Y,g����D�>�w�,�X��㑠ѷxv˴W{P���*�M�W�OC�N���<�@$oZ[
r������|ch�����T�(A��5�/ÿ��-���-j/�f2k�DG�-��%=�|9c��Ք��R�`&`����+��`�ڎ��c�ٮ������5�(Yx�k#����i����AdE�܏���F"�Et�5���JP�,'0E@U�1ψ�����i������>X������O�a	9�tiS�')���@;�;��)Rя�is��*3OG��n��.aeL.�P1o�lar�����:bM(��o�(q�m�/�=5v����������g�#�QafE�Rw�
7VU��}sL��Y�Ps<8�ҽ���J��qad�g����:Ɇ��d{�pӏm�N��tqw:
��eб��c뢘�a�R�ǝ�ݼ���g{e�Q��Q��!� �(~9�m��F'h��?�e����857�����"��v�s(@�F���Թ��]��d�LHa4w�sv�C�C
Ӛ�<z�?/���_^Wc)t�K��^���x�����	/��e�e���:���b���&]�)t-�Bx��q��h�?$oޠ�鍺�>�*�Rˉ�ߡ K	�b�QV��C�V܁`�u'�;�Ȣ��0�t���	O� �9~	3����-۩
�Q���V˙s��7홪�ak���x2}�yO��2��)��a��t��pG�ޑ��k�~�a�S�$���n � ��<�M}�%F���4J�S�Zk(C[�;v1ߙ�hn�a��Y�i� ieK[��Imm��L���� �|.���si\�|�?:O[Q���8��3��V��%�Zϥպ���-����*�w�^]�ty%9Sø�
My�_{W=o�c��M�׬�6� ��d�V�J�*J��pj�Pq��ݡ�q&�r�D��͂��S6\53��N|"�_�^�͕�3�G]�z���O%�k�m
���a���%J���0�-��01y�j�ώgA���ћ.}�Ol"!ߨ��ȋ�W��k����a|��pC�"j����P��٪ԍ���n�"w��>��q>J�Nd'l�̯ b��@/��C�����Z�It��
q�I��b��E��)��`B�K
�Zc^5T��|��dU��-[�C�"=��so6₩�|<��x��n���m�1*�uX]�#~޾��q0�x�3"=I=�#�ZC]����E�C"�cDy �\Q���% %W������������ȥ@XD�*��<$O\�0|�0�W�_�ϪWr�tߟ�||6,z�?=�����w�.�μ"�yG8�'�5�lgy��Ά�U��zAB2<����Z"жF����-��m�Ԛ�l�h ?�9)�{�%ģʬwT���d��v��Z�����l�)��ryQ�"�Άe��ȷeuE�ʉ���I����K�)elѬ)@��ϕ
��G��G-��'�˵ub�����O��>~�[�������RB�b�\�}����uU��(I�_����/�	�Iў�� �Hz(�0�k	���1��X���ƙ�Ki��zޭ��Zdn��=v�;Y�S Q{_;�S7~C��+���y���J=���"늸�'�*��n���O'| ��sh�D�2��ݶOh�fx�WJ?+���ؘ"VR��3�6��n�&��!��i4��W��-M��ՆOç�]<FE�*E�pre2���M�rJ��n]�t��2|��c�(h@q��)3͞ǘ�&��붓�@�-�Y{)zN��[�� �l�ޯ�z��Ȁ;1��Q����7���n�g�'�A�BP���s�;I0�_���}-�Ԅ]�8��CI�n����J����C�y�i�w�h��u�����L{�3�)��I�ڊ��
��w��h{�m���]�4ĢW��+��:30��5�X��=&S��y�U���$��+���k�,�����62[9�v�}��e�n���������T����_��E����K���}yV�$o���P�x��Xi|� �ʷ��q�7*�/�4
�����ks7A����¼@��a�,T�_6��7��_�,z%�����t��h�mA������#�ծ��>R��>+ڃi>��u��8�6�p҂vA^�	���� �İU���۪�ǥ����������#��m�ĵ�đ��'�o��-�K6V�oQ}�u��ъ��`=wJ :��0@r��%m2?>�;��׃��D}E���fgJ��yO%ҭ��ț��JXE�#l:��/��z��Ǽ��t)0�bu��m��'O�I�)6Qy����M�99�Ak*jY������ąD�U[�Ī*�:{�����5;��&<��ԧ�<?(Q��[g�٭�eq������������k�n�,c��aL��š��s�ՍW*z���\�0o�z����ujgR�Ȁ�_���8SF�A~ȟ;�x�ތ�x�.vb�_d4$/�s�L��&2�
�՘�C�c>�~����Y��o��h��D�^��`._�L����G��do�z#1�|�W_�R�ة/��kz$e��kZ鹾������+&�<���#!�P�IC��M��
8��UF2���s�﷨��Q)����������m+|�	���&������Ndz�s��.��tW��5WS(�3f�.^���T�ܶ(Z�Hjf��8�8D�HN*����Nc�3l[1}g��9嵹,j1�ԗ�+��&����o!��b�'g�!�b0��?�}AW����$6��5n�盋y+c�Gx��֒���3c�9��u�w=s-lGM���� �T�s-�?���������v���;�%����J���L��
s�o�?�1��bBlU�^�.�eFC`�=�q3@�+j�V�͓*���*c�/6�l�z�Yl?S�YdZٟ��4�1�[U{>�,��t�kiȦ��7v3Q��emҎ,���"SY�A=�]RS�ؽ����%ʾ�$����$C��벜Nh�?���)=��KBiC2����M�ď��K����*<м�������M\8��|һ�ݨQ�Flt2.t�Ii����ܡ_�>���7;�`5��V�Ge� Ō���j\R��/��r�����;���T�n��ŭ	B�1�KLs�m�{/��tq[nB��G����KM�_w���+{$*��6�O�đ-���-���X�c��g���ȣ��]Q��#
���u!B�l�HU5�T���q鼈���ö1tG��Յ�ӱ�q����X�2(����?k�� ���<t ��mwÖI��}��!�{w��V$ǔ$�~��t#�۬�M�Wͅ[��Hl�y�ɤ���]ȦG�)B^}& ,yez�'
bfҋ������&�cv>��V�����@(1=/�8���lKK�WڨR���I�T�X���7�qV�w?Yx�^��� ��s���5{�����s��O���A2�����vY�A���UW���
\6h'����3��(>��E�[.���s3��������
�B������O}�")E I�6ۘ��~hP�\ΪNӠ��ɉ����.!�5>6�Y�;2�O�	W����YT��h�h�.�"�7��Z7M����^�ڥ�OR�d����H�W��Л7 E��/�t�����n�q����i_�$`Ƚ���]�o��p��7>�D����"�!�s>LVC,���'���B��Q����o�� ���&ڈ���:H�����v��~Zeˀ�XbvC�/�UK��p����*s��қ����R�:T�&�
P����;�R�gɘ�Od��M��T�'v�-+x�h~��$��or�o������
����DB)x��Y�
yV���BW�<?G�Jr����3`8�_R.@*����6 �?�Bק��E]k,2�5Y�3��}轢(�b�S`r�QP����*f�,������2�W�󇄀NKW� }}m�9�0�p'����F�Fb��X��$O7��SV�>]eO��}���Amc�FX��Cխ8[v�)0t7���9w��;����r���K��]���7\n��ŗuޫN�?K�a�v���:���>��NZ�On8����/b�6@9��k������G=ߝ�)���J�6�'m�*��[�xh\H^Z��_��'l,c�2S��/��.ᤛ!6	 w<� ��Ȫ�*;�nפ3��OJK�s@$��dt�q`��x�0���AU��k�z���I�����[(͒C���4��F@�����:yɔ����@z� ����q))�ǩ��h��N�yB�@�0�޸Zȍ�K��A��6%*��=G��<�ś����Q7?�H�
r}�w�M{|͌?�H奵!�.��ږ��l���kّ�hwݿ$�6/�'0�C�PM�{[�f�^�8�
����=_��!;F��(�W~̾�k��Aâ���,D�^�Z+�b�3���~���k�6�a��&�=|�PC7�����7N���x��	V�)+���W���=��S�I{�#��ɿ�gmh"f, ��+�E�Öx[r����4\����*MA��] ��L�F*��,/�Đn����&�fO&t�݆� *[/U�6�&���p��є�)3������Sq�1����bӭ=y}�e��y�-�.yd
����iˉ�}��
���"So�+��~R#��O	벗^v��%��W)��ǜ��Zߡ�V����P�6s����%m�Њ���f�D<c�G��hߔ,�gb��K[�2��a����T��6��X��m�k�΁_�ř��w3����������-##����%�ڑ=�k_��{m"zK2��r�k��l�e�a&���{/)�K���������z����Rn�u�-��.�&K�@]�̍iH۽d�fH��]�΍	R�R����<��ĭ�D�k
�+]����KyqWgds0�Y�.��C������sH<���dV�~��|l'tQ=�Q�'|�i�aQ,��e�1�|ꉄ��*yC�a}����q�~ힻF	�6��&�k>N��]O�p%ϸ��N�c���f!4B�q��v>$'�����][K�R
���+Ċ���w]��%,�*#��P�֚��|�/�'�Q1slP=�u�����Xl�Ձ��s��@�m�"����Q�^Q�t�ۓ���8��o޷?�G��-�9x����eˢ�����ŋ�J����8����������v0������T�*_�KqNu�*�����bO�;�8en�P�K+�8E�0�T2���b��"�o�Oe�}�!�5�O,����H���Q%���ɷD�w�_P����[:ӌ�-�)UH�׃ ���:Խ��L��Ty|�8�� %�a� ��B7{"���"�w!�3q|�oD&%�}QHT���9�1��m����6�X���Zo�j���;D.NI˭��Fct[X>�7�N��^
F�dp��J�)��c�t��["vڿ��J���F\�H�-Y
��|��D*�0k�{�l�	���0���*p�iՒ 3���o�`�]�z.�v಄������]���ޏ�q<�S�iʌ[�d�E���g�Q>�%��r/�4�z�^N���"�w����b�.*������)�jB,���U/+�]V&���j/��2+���Z�,E�H��f����Z�fä@[�\XOxػ��F�';m/r���.�'￘=~oV��9͹}��k�~�w�{�Dع��� lH��(�
ݡч�t\�o��V��Θ�� -=�w�򑰔�ȕR!��I&b�d
���M;����p��px؉����\ػT�V>\�c؞Ң��\)D�ɪ=G��z�Y��;O��ff�g:�+��,��-��?���:/ܗ�O�ٺ�7�ޝ<g8"����=��|�ݣ{����ۆ�́����m��eij^��;�NO8��{��Rg���߲	6Mz�r9*z���9HJ|�3p�t���\�ͬ�^h�K�Q.NP �4��서�����Ǜ�C������W��B:#P�)|ޢ�-�{�J�BNI@�ק�8(:#�V�dsm�8*���хd5��\Tt�#/����\a���e�n�9���'ud�~U'��W�p�p�p��4)�R��Sn���$�HSb-�.4���i΀� ;���5PE�=�e�D��B�G����sE�7�1�z!8��}۰w��w��d��y
��M�g�P�K��P��h�7�8�^Õ����u-��I��e�%���-A�$6H�j�?l0i%6���z�ʐ����^.���FW�=-'jE�fv���X���/ <JZ��,���Bo5a�f��(���d��\8`)8d�ī���K�m�k��,���N��'���꣍�Kt�_��xr����u���|o#��/U�WbӋ� ���6�Mu����k>��T�Vh��T�wV����^����ќ��K��CI�{����A���2�/�ȶ����z͌��X�+�
�-���8k��al�v�|�Ea�&��l��;?V�8v:0�c��x[�6�Ԥ�2��X����Y��o��q��5,\x~y�����
*���1�U���U2����-��]v��R�t��\ �k��K�HD����ͭ���^�<'?�c펅�30/N,� �Q�s�旄�7�{��X�4�Kg
s�"�KB�dj(�2�u��s �?BOI^p�!O;�yU���i�jWx����J�8�L"�e�Fr�g��JIi;6�)B��w�;5�X0��x�x�U[a�W���� 5�ARތ$x�V4����6�Q���W�٩sW!������緞-.����)��K���8m�p��v�T��_I��� )��:͇t�W>��;2�5z^��Ptr�2�\rwr[p�$�6��������L�fK;F�rXP_�z�L��Z?	,�m�N�G/U����/`�G!��/�s
G(/�"�.5�������F���A����E���
F�8w�焩��[[��E�p�68�^
&d���R��L�3��Y�摼!��uC�Oo�s_[������#,4� �z7�,�D�]�G'�95$���w�����uV��~�D{7��!�dR6����,�'���%����=��񐏠�:i�wfA��彸���<�/�n�ŎoҤi$KܟvF;���DG>L��b� ���+DL<��ũێ��ƨ��
j�LDr�b��h(���M���X�f�=������'Br���c�_h�nŝ�lݶ�2]������_��5]b*��:Wqh��B�zLa��`ۚ���(�����+=�9������
bbz������H���QR���T�AM�L���uI�M�����3sߨ����Z���9d�S��~M��DbIk��>��g�6R�G�n(6ũ�\�;A�0�R��х�v�Ik�dW��Z�˿� !����)"m;Y4���:I"��t�	���rm5=�}S�sԥ���48�Ǹ�f2�v����mMG�=��9x��Oen#9?�T�8�aI!���wK�k��nL��~[I=�t#Q��g�&Z�����cJ=�,C[9�O�j1��0�>���N����l���e�������G�x{J�}m�����0�EEBY[ݔD2`�)1c �p��S1_��_}5{1f
��V1�bU��>�mm�l���\$��u���ɠ�2��`FW�+�8L��l��'F�WI����o��C���T�hE���uo�o#<+.�/镸�/K�;RB+.q�N���[�ٖˊ*E�3�JP~�ެ���[>�(̻��١j�y���j�$�����k�OD�2��K�����P	���e'�Dp�U�Ø�3NVMb�E���j�d:V��P���f�KըARW�HՕ�%lx�S�w�[����u�P��B��Ŭ)�(lҾ�j�P5��ek	��3{Ě�)�8ߎ� ⢔H_�|L�]�y��|�235	Dq�����B�!��4�6cW=��Z(�[q2���/[�M�ӹ�BI��2�ыWM.n���r]��f�Wr�*7.��v7O�x��e��EdQo�]=��VJ3�4Xy>�ܫտ�j��M"�����s���]�L��DيXrO�	${�Hq��A�=�d�Ϙ���}h�ޢ*�*R���8��x�#���>I	������|�vt�b3��f6��R�+��:*8N�i�'}!���AXxN�g?w��ݾ��5�?ҥc��!�Ԏ�p��^���}Z�DD1@e� ����)8 *�R>J��ja��H�!��`���Sl��&GNDT�R��#N��Oa��Ȫv��tN�y��mk�e�rt�SGU�Ă#Tw�v+t"\E9�[��	�|*�0���3�v������E {)��O�D|������"
	e����~�N�5F�)F��N�j��ۥ�(��@ۅ�������6�P�c ���Ee�跰>�;�e�}�t����y��L��7R�2��ZG����XC%����gC}H.���n_f����$�Xl0gQ%y�߻�d��!i��c�(z$j��1���[4nM�p%_R�[����{�*0t\�H1�&�X��Åz����n��C<B!�=���n�/ʜڞZ@n|X*��4�5��F$����z��YKv4ϿO�k��1�m �ޗC�ʄ�u�ɶ\��L^�;�v`���sV�)������i�h��|m���J�+�"�8�Ζ���x��^�t��l_H|��qH�=�[�����(�\<yd���,�;�Nw��l�r���^����.Vm$�i"�(�6 �ނjru�x���{�q��D[f�w�\��� V~_��V�
�H�r�ޏ[%�P�3)&D�]a<<W�'��kM_%X��>����>]�8���A&��R�l"�{��A�;IJz ���&)p�`��4{�W��\.	��ҩ�~�*�t���u�M��xg��NO��%�}kk��>����_{����ϑmݥ =G�bݕ�CԍhЫb�M���1��H b�|�/�z��r2����$�e�����f�z�݊}�Gc�l�/ͦ��G�����
�d�|g'�4�<��ϳ1V�G�� aKҩ����6L��;u8ms�@WY/����;��l���C`��r���h}5<�2/��_��_������wUk��X^��mK{�*���k싎�剡^�&�ICt��I�����6�E�nE��iT-e�B�벎�Q��Q�hsԬ����P
�Z�{�������#
�zp�G�s�����8�Բ�yku�ynO|��aGs�Fl�B���8�O_̭k?�&���i�.ފ�e�}����ݸnC9��9�-��~v�����G�d���D�w�ZE�?^���m��������6#J ��Y���R.+��~}���?����Q�a�+02�SJ��ad����7���z�
�1�Y&�?{]L9��=�?�~j��z�c�I��a2�6y|�+�JlH� |p��a�[txp�(�t����\����p蒌Ӝ&�y��#B�wĻ٬�g�%�LO�P�&�Gآq��#��8z�ì#���9���bY����摕�5������S��0��%$�ڱ�_=X�yu�Z �v���d�PZ�7���x�य��&g�șwa��` ���}��4���w��u_(�y�yȒ}���W�O�����K|Ytﰻ�EQq�^��q����w�-���S~��3.�v��dUa�]�g���7,!�X��JP�ӕHe��ڋ�M��s��}���ɍw,��׌˽KN�.o��+f �*(�b�y�G%Gv�#Õ���!�����$�`5m^AnT����.0.թ�W���j�2�b;$&��( � �s�~��3�F�;�ȳ^��|��?��<&N�yR���~#���`�1&��B����%k����Ô�.t�zh��J�F�YJ�[�dl���v�i���ao�k
N����MF�O�i"#��p3���o��>+��&-.dr��G���FCۺ���HyYuk�d�K�$�i�vE���p�j�^6����I����i�bv����ZU��|��*@]L=f#��9{���F���TR�VDi~�A[D��	N_hOo�-)�1�~4�5H(a@!�!�2yA@Hl��J1�y~�A�cb_�.8c �L�MbCg�T�8�hb����bN5��|�~�\Zޭ$G���Ge�4�sn���c��T��E̳q��e��I��f�C�Ԭ�޸�Nw�iM�y��8M6��3��5v1�#pV��m����)�b����8�I�>��O�Ydx����'�&��\
>�c��Mɚ$5��E�*>�:�'��w�:@�� �PXw�`$E�WаWo�饁��L�!��>u7XĴ@����Q}��1�����Į��J�'��7���jAs>��g�f��h�ׅF`Cš�{�u$F�#��T�.QP�'	��<9[�g�i�����V��v�[�G�����%��F�8 U��_���F�I���5�<�j�o�M�O_�T����ʓ潳n���x��A��o����"Nk��#������}�L��/���=�FY�XרЎ��5�3c,����+��V~�N5�)L�8��0H'K+��xVp�qw�m����1�r�v(�m���WE��g�ao)�	��#.d^%T�n��;�$EW�ïe6UĒj;�)"����D/KY��c�[V�<+ᑨ=u�S��Ԃ�U]�?I��GU�j|��G�-*��χ4&����a�;�)�7[��i�
"ˢÞ�R�w\��Iʙ��6وDJT��h�/�=�9��wH1xBy�\��_��tWfmS�ܝ��|yIu��cWsZ�ZI�u�j�ͪ����{��k��S=aʄ����F��B�:���j(���������y*;�>�*�;�g0��)�r9����>�CvH�;�K[��b�#Q���"�����BӨ����\�pOL���뜁ĀGmL�Q ���"�-����,��U�o� ���
T���ʤ�nI�^l����
FZ���?�����1kvb�i���j9�7��1������"�W�^h/-p�.������t�j�;!�K2i`�0|,��cz���p�4�5䕹`TN�QW�I�.z�̘����KE�m��E6��vf O 8Hl$�X'�9��wb�����m,���8����cf��SXR���.���{�R��x������k��)���b4Rn�/B2�P����в��L��l��a۾鍺j��ʆ�` +���]�j�*5�y	�)������ه:h�2��dF�i��'T�����B�g���1�ذ��uL�7ܽE��)�w����#��,!�|�B}ΤUN�XqC��2>�NR�t���;Ɉ���%��46���쯨K��?{���`v�p�>��\�����)�g��$�¨w����V9>7�]C[Ó��G �l�����O���{�y�<-�d�~~�j��UԔ
z>d�4B;�E<�(���7�gŢ�Gu�wI���kEG؃(��,�],���լ����	T���+)]ƺ��W�א��T�����ݩ��4�{tɺ��9��b��z�@a`=�.R;%A�\$�|�p8���F0��Z�*W����~�Ⴎe�n�Q�[�U�zR��/�P*/:)z��Z��ќ�����JvxM�2_qr���n�� 9��.u�S��W�Yo��;ݟ��sp�윊鿑�y�*>"
��ǅĄ��B`
�wJ܈�����X!��'��С�
	���֬�EʌѺ���*V�0v���b-�����OA]�Z苷xu�����q���R&WqMѻęV�T���7�v/��*Ѭ�F���H#�N�9N�{�e�m�M����DV�W4�߀�Ļ�k�Bp�0T�+(>I�Y�
϶V�.Xc����y7�k��/zY�r��L���}a����I���l�̯�7�P��G���=5\TeCh8�W7gj��
q5�yy�\T��+ܯ�Z�3Ԡd��ș�,ڷ�Q_	l)�%�?ډe:�%��\I�YX/��T*���T@���u��jT��cX�I*�F;XH�0��k����r�����BJ�Y�N�\�X��*QQߪ�J��Ê}�gr��q� �<{s��+���,��!�9���R�)i�O�E2�gρ}P��pb�������Ȯ�H�e�t/{z��e��aA_�mh��]��,E��H�P7�ݶ�V��۰�����!�?j]�?�:x�ju %�k=n�Nv٥F����մP/��u��!Յs�黭ҋ	�Z��]UW;�a:q(Ǭ�P�c�k�_9�:�CkF�pU��p��b�V�fՐ�˸�Q,ɉ�Ļ��!)~W^2��w.r;DV ��)̷}Ӥ8a|�9ׯ.C4��/���(�쵍�@W�d`�p<=3RO�n�bJ�C^��r㳠M'�6� !Q:�j��*�!�úE2S���i��R��ɦ�d`�=`�E�KTFf>*9��f��4D)�`�V��+�P(���C�����u'��5t?ŀ=F��KHv�����`mJGa�#(-��0�}�e�8v�1p�|R�b_'ơ\6�ߠ�$G�'�ldqr0�j��P�N�Ç�U�H8 �=U|e�Z�6�t��1���.%�[�P�.p�B�0y��:��m��\��|���[GY��l��[;l��,�8k�;Y��{�K�ZH�oÇNN����<���r裐�펝Wݡ$�M58j�ky������w�.�;Ab��^bx��Z��)fx��"��NU�6���
��PԪ���m�y�V%{��p�0��q��g6�go�n�a�YҢmں�w/#'��w��\�8��f��Nn̚���}�{���3�*�������y����A&}_�@
}�]�.�IUܜnK%ku:����|����`�[�;'k��$�����ܾ�����f�t�H"�P���f���NQ��py��+ע���:-��	k�Nt�X�0���N++�H�R��03�T�I���_�+q�"�9��&M�sQ��4ӹ@�W;l����8��X�+K�}���8d��7kH'd�Ν�Q3��!z)C^FU���xєz�ݚ���ԟr����ua�=�Ќp+V��6�4��gR,�$��!i��<��Gd�)��O��
�ڰ��=&��C���\~֢��Ji���L5�֟��|�?LQ3Zq�8=�>{"a�)�M����қ5�R�i�}Ip�D����g�����R�~8�+E*Pv�i��v,��tv�V7��J�B�y�/"��+&�r���u�6�J���w��8�;�&�4�N�=l��!C�ձ�`�ة=��b�Q��ϷI�a������E�� PU{���2���C*G#b��VD�Aɝ	;����$?��.�XR�Ѓ�N>N�:fH*�ʁ�YTjQ����y/F�^9��-�	��!�P�ݗ|��u�!��㵅���,U�:�O�jhZA�7Z�����X�9'��tʵ��mݣ|��;�'��Y�;��D�ײ�~=��;P}��gG;��Y/��HU� &�2	^��FUj�;-��ǉQ���a�>��b�|�Ji1��E��σ�x�~>9~�s�tP$�I�� Q;G����������]"�\N���������KL�-��6x��Q�H���,.KU�U�'�F{��é���s�1���Ҁ�7�x�?Jp<~��x����a�z� ��.����2�^��yMT�ю�\�����$毎٩է�c���
�W�j&U,ݑ^���)��~�Zؖ)O���x&a�7�e%�p@n�-�^���U����ON jx�����ܱ�z;	�g��_K!�36���ފ��/�>&2K���/O\�e+�uʪ���b���mإ�xYtAS����藎7��>�~��x�3��yT�pn�лR�<�4�c����˫�����-���3��LI�%m�&�v�6��c}���«'�5����)��7���;��,�����c��>daH�';4*}�^4Y�����7y�uSK���+�$T��ж�׿�~�d��j߻��dף��/?y�HUN�����j��Q6)����w[F��XR�_E\R�ث[��%+���7R���p<�S��]������2��eO}�8*��0a���h?�f��[��+�$С��P޽�ji�@ �[��\�-[�B2�A�C�1LI=�|��[8��[���@�[_sE�@(��X�J4����a�=F��I��n�p<z_�J/��/F�.(��y,��J�\��j%��k�l:�k:���Ɣ7S ���=}طb���ҩ�*����y��5�{Sw����EET��ҋ}HCQIBAUg�Z-�L�SQ:�����bJ/
C����
�d�'�0���;<�5���+��K�O�Y�=ꏫK�FTa{
�ܶ;o_��U\��f�d��5�Q�Q��8��/�
�0 y��l���SY��D ��/6��Q �#oFXs�?[�R��.��J��Xf'�V��ܜd^����2)��]_�9^�J����D�RA�m����ܡ�׭��4Li4.�3�����"��o�'c���v��~�5B-�)���g�b�X��-���l`g'M;LN���`cgSQG�j
���e��p:�?�e� ݗ���؄�Z�@JK+��kx���B��=��P��&�z�.�u�[
&�����������$Z��P�p��`HI�t~��\J���g+�1*ܴ$�H3p�,|�mQ�I��t��`-=�c�O���(�z7J�û!oA������<�8��j./�9�u�`ç��lnz�r v:�˻@ʪ���ބ�X{��K�k�2 f�Yz���������N�it~Ů$�N�s}H<*���	���g��EW{Za�&�H��I}.�<��i��1��@[��x,rȊ�Y�r��7�:�
�$�~
h���}�/�w�Q�%q���<�2���\F�{���%��.�C�h��@��0�>Z�+������Q@�:K/��g��m]q��u*�І�4'gR]�����\fp��Y��ce>FOi��?n:�r�%�۰ ��Y�n1kw�~'H�����]���s�|]���5j̛���GԼ�#�us�w���8�f�h����
������4��y���4eC��K�/xE���>��8F�>l��l:�_H��g�Ι��������Y��7�Mi�O;�i��[H~�l��*�<�z]���(9���=�2���|){-WyP/FMzW�;=u�mAq���Ѹ���؄z���1��?���TIij�`�E1����~���Z�܊zYQR_���AY��T���Q`ײNT�~<�>qSS|2��G�#3G]bC"����5�ɻ��4|�%?�#�$��]������&��+z�#�v�r�7R������y�>���;���bĞm�{�� ��ac6A�獐�f��:x K7�r���p�VT&�#dנ\W����q��|/�<�I�T>�P�� ��G�P��OI�������d�:-{Ӗ��ͮo穰�6P7�mE���l���HkI��ћǇ��u�]�K?�TK�(8��xr�j<p��4�Bu�H���h��s�7�C�PM\=�|����~{Ih�$�@�R��S�A�9m���}D�m��k� բ	5!�{��":/�3�(����3� �oh��?�oqq)*�:y?9�������Kn��̙��n��ۙ��8�$hw�* Kݵ �~���G��4��#rh#�ML�2V�$�䘂		þ���w�2�y������|'�nxrH��ޱ�ql�H�(�!rY����,yc��n�?�.�yg ��V�� V�dB�"���!�*қS ���jPM�;a�OuJ�|�1�C�<����� &[ ���j-��fґ�])�K��/N���[ \�Qq�g7�m�踫��z.iZ�cH���HdI#����<Ҿ&�,v�ynKk'ڢ<ٽ�p��s�{\D���N=�2%�"Q���d_�����:	m}�^��G�,��1�-j%���8�W#Lp����=�Y`] �J��+�C�{��o�k}lT2�x�3𗰳���Y~#�M�kA�E$]͙pW%��d/|�L\���Ψ�ҁQ#:����U�K�V".ux��NqUWit_^}�����`ܦc.���F�\�E���7Ņ��4?��ԣ�����k(�G����\)%G:�8� Qm0�P\��o����9^E�A*�h5����7coBJX:��D����� ����D�vW2ڰ%�|t}���H��S������g'M��p��8f#e:�;�k(w$�Z]�?��R��/�%��&�v�CK�+�/=tHf������ύ���;�~�RR�8c��~tKX�3m�?h�}Jt����u���b����	��o�Ҩ�n�^�!4l�C��k�3 +΀U7#Ftᡝ�ǔ,8�푕[�+@1�vu͜��W�#��e��	Vs� ��۶٠ԍA�}�NI����[it�(�8e�c�.���	4�K�MQ���F�˺c1���f�?�O /���m3"�Gt�;�,��G}5�N�[�ތ��cx�,Z�c�Y�}k��(��-�	����y����.N��4C`q�'�!�Hl�9�<�$��p���W�k4���ԋ��k*Y�c|O���t��G�h�5��� ��}'X���Z�������3�C�F=t9��chK��[��*�e���X~+�d�RCIeYt��T����U�?[m�q���h��<4�P����@� g����ޕ�^N\R���:!�d}��s�����2s�u�6-hsՍ�-k���aC��vw��l��sE�A�h���Fx��e@ֲY;n�P�Bg�Y���Mv2�f�l��m�M:p(�	G1����t��8O�y'1y���'��{��H���+	�v��$��l��`�%G�1�N%CO�Vn�^�Q��<k��`�a"s�%GgC�2�8oO��7��Wi#��[Ѓ��Ģ��)�4 x~���Q�}�H����DP*z��;��g0���4��1^�nu�Zp���Rm������/�5�bmM��-{`�c�u-���b��������ٖ�d�l%���r'K���ǵ�\��d�_��C�� ��̆Ҵ�9�Az�ױ�(�|���#��NꆠS�T<��[�z�`��� ����{�س��҅�fO>+�)++��>uZk_����,+B�adq�T��x�+��[}Q�iPa�S��q������13��>�J�0[���I#���O�_�r�ơT��]Ҡ���Ty��:A�OT/)���XJ�s5]�R�m/T�\e�3�U�і�Xvb�Tʤ��i�:�g|TX�_�RԚ�Լ��x*A�8ͭ��B�1��,�v�R���X�����^��Y�q�h �ö����j���Z���P��e��폚�'\q�M�y;Y������.��h�a߾��a�q���F�`��x���Q9Ɖ|�$.-�����^�:�K�OV���75�l�l.Z�*"�w��������#����G��BF8x|�s��hL����{ű��u�>�GWJ?��Rۖd�3L+'���,��K�y����h�moX���j���*����b�a�����Nq�fb:*�k�6�C�Va�T�	������f`��=��q�����C!��3�2ʢdk�/���W��.-(��="��z�L�K�FWVDw�����\�z��o{���#B�溕�g��kx!��������qd+�	U���V��j�W6|�Ώ �G��@�.�,Z�t�v.R;���Ү����'f,�����I=S��4��[6��|!�t�ɳ�,T"�)ڽ���
�84f�q�ݗb_�[�S��[
��%I�eS)�N��i��Wp���.���x+euu��I�G��@��%G!E�8x���IO�(�l_�&{C\�-lW]���,�� A*R(�}�Y9H` ��C�IveC�g�]��Rm���H�OT��T�>�B�K<׬?�;l�Iq^O<���5�7�p&B6;���a��c�:�ѐ W¸�H�7lH�mt�4��fn��5B�͂XrH�|�Z�џ�yS$37��RŲR��^Eo��cRK����$�$��yjXZ��hK��K�)��+�F�����c��M���:�ͬ�Zo�M;�猡���βhZ�H��9���aT�~!�;��_�~��)e�97�ח�e�W_������n�����Y.w,�]�h�i��c��-�D�sn�v+���͈��3}�e��3�m�J����[������B!����W�p��W�|���{rY��8��WpE�;�n�{W��T5I����"��|�k<��L�"(9YPୱ��R��Ɓ��s�����/u�/�2��n�k����	�+� �rv%���|�z��Y��
�+�h�hg|V?E�Z�AW�y�&��Q���8��5u�9�R��	�Wʦ���/e��o�tg�:�7
����1�i�_H��[K#��F�O���~����g��B�˿���*���n�W��?���*fe�k���u+�>s�p\G����I}�l�{����ұTU���E��m[d���}�t�? �7(i
�	u�y��N�w,OYy�B@Swv�[���|fٝn�
8��q�q�R���e�s���+O|�F<oc��ܸ�	>5����$
�N{�Sv��Y}�4ܔ�������R�?Ѓ?!L{�����(Vݜ��>�"��u�;%�#��~���F{�P6�������@�+��^��u71ppBI�Ṛ;�����6�&�E�v�0���ُ�ÿ�t�ּ�����C5/���n>+=��!rh���\�v��t`�jc�򶧯�z��9��gw'�V��!	��ϭ��c�����vzߋ�y�3�9��'�*�M>`�g��{����M��0��ד��v��)J�'G�dDp�r�h��e��r�Ԩ�����Lu��xd�(���Mۤ���eVJ�MzR�|g�b�Eې�G����il$���zZ2*�ը�+_�@cy�� �a��s��\�l�����#��ygH��LM�I���}�A/���ŕ1�V��S�����B��
��+�/�
@�
^�x��f��ޕO�Pb0�]P&B4�{d��S�^㞷�4�E�p��Q����b�T�"O���b�-�.���WQ��x%O8�_g<7�*�@ڬ���b�)m������ǋf���Ć�ѢCg�������w/�9K��)8
�g����=[uY�c�W��� �F"Jc=����Qǅ��'�g��8}���ݹ-P��P�#����X� ��sE��%83#�/7���s�D�9	G�F�,��_Xg���K���j�����n�BIaSYvf���~yG��P]Ie����\u�Ş�
�
p>�z���U�';D��r��?�p�͸��+��G�k���E@�K�H��`چ�Qh9���<�9�<���
=��(q(�|�8T�K�/���[��VO���(~r��Ӆ�r�l��8���Q쪼�I��,����zxޏ'��۞�9�:������۹�*q�B�p���|=HM�SI_ԌpA�p�GT��+A��6��\�a�1]U&�2����_q�'	�Y���"�Uc#�J��S^�6-�2�^����V�,�:8 8-�<e����3�{��$E�˷6�S��d�Ԛ^k�[̦��;�Ny-7�2�Iby�Wlr���CA��κV_t�Ji毁!�2��7�nY*d"C��Ե��(0��GS����p�ۀʑ�����xc���m.�NDyp���.J��!מ��~����a5_��38��<5'Ay3��	�|�m����𢁔${��%�r�"��ٹ�w5R���Qԥg�%���?���8���z��τ�j�^P�=���'xn.K�8><S�0�������*�Ԝ?(r�\zQqحB�k����Ca�L+�9��1lj�m�^�{�A{R�Y�n� eڕ;��#�F�*ڬ;,�y�N�c,����QM�lf��gk�_�q�?��M3륨��z)�k ��Ԩ��*12\�#X�3d�!�Is6��i�Yy�.d��)k�H�Ebr!��݂�� �\u�ǰO��mU�W�T�?��AC_E�	�uE�;��U���gn�au����������vh"{۸��'���S���?�\��C�@��x/�o��=?���*�D�4JU�O��t%��� ���G�BIv���!O��pc��W6&A�n)���-t�d~��c������:Y9�g���%V��S��i�@�>��Bc�r@d8� ���r�>[�}I�P�g����'q�3���kj)�F� G.�n������=����x�<#{l�4F�p�.�L���c�ݦ޶6�UL,��C� ��,��wL��Z��E|`�43����}���oD$���j��������yuC��=���̋��0�7�t���G���Ձ��WF)���^�	�rM)��Z ӅK�[�C�z��]�T
G�p.p�l~_㛣����O��ɮM��t��p<�K�֔k�I2�h��P�=����E�[�u�H�.W9��_^�2|�w~���n����6�*"���z�]���lȓs�����h$�i���<���tovm5�vV��R�0��F�,�[AX�Z�:����R6��q*�o0B�������Ԥ�t����&�q9��>�Ϙr������� ���������d<��.�k��E��I�����R4M1U��QZ������.T��!��0��i��tt����עu�2!���RB	�G!�e9UG�C�V��g#�K�N�Sc����`CE�0h�z~�z�E�ا�N}Рļ����c0�<���1L���T�j����?�*p�8@0�X:|v��._HƟYh�l6T߯���%�1������73������r��j;��p2�)�%q�a�W>��. Y���(����GH�,1n����9�� $@ۿ�
����v4d�¡1ڭK�� uS���ޫ7L��P��g-)��2��K���-���2����5<qCA8���RҦΠ	��VD%U��5y��2ZJ2��]�E.�r�B0p[z3��Я�V24k����EJxZ%8��� Y��6rǛ;�� yj��F,d��
����q�4�47-�� D�ݶX�r�ly1�����W5T̝��7���H�g�y��k�3�� _La���H<eJ��9��l�����Q��v��m3�m�NF*J��D�k%'W��G�w
�� 2Kt�q�_���!ɪ��yH���O��jH+���"��QY��r���r�l��S*������z1��Y�;��TR�Ȏ[�2��KFZF��W�䘹��Q�4��.B�#16P��@�7����ȾSJ,�4������;�y�b���ơ e6/G�Q�z&;c�����xdȲ�VO�M��kI��H!��G��6N�=22���ˍl���rb�s@��Y��8l͹��5]���X+y4���%u6�Pc5��.3,�l�8*���ٌ��,�RM��4N�R��T-O�#�-��m�1�o'Ȏ�qu#�r�������5U�R�|M�錣I��NS�%%<�eɷǭ��̩�ޒ�&Z���L(��c�5E��p��+3Ǝ"Jn�6+�m��|����I�V��*f�t���,�B�pH���X5l���	�2�X�ω���,g�$�֔p���l�uy��B�	E�}1��_z��%�?���4Z�<������[�7ݓb�.�L��7ťDh��jO��E��(7VK+|��he�hEj�HgfNKE!�T�J2�
"�<��&2Li�hqHzdRL��+f�G�
0��y#R%�J2+l���ȩc9Kb�Ak+C�㘹��S*W�;�Kʾ0�����w,Ō���\��ъWچX��uǭ~�q:7�Ҽ��5ىt>�ɍ:�.���1�野Li,�!�q�/�|,�����1_~VjE1<p�������FFfR�c� # <�E@���<-�8��u�z2xq 6E��&�e/���:����&�Xș+ə-Km�ab��c��Q]�<��_���͋�ޘ����ni1;*:�&��u���V��WS� N{ML)}�uc.�-yb���hȲ�*S
y-�1�ͪ�G�Hp��nD�����#�c\�l��)�������,�A��Q�
yŌ-�D�,
 �9��U�#���%O�#��q^���p�ll���&է�̞M1U�u�&8�y
�3܄(T�yzc*�Q���k˖�hB�*=�[(ea�Y�x�P���0��:+Kt�T�[�DL�ȹ	<���~��(��`_f.P�c��qH�e�s�Y�At\)�x��3Jc!��7jL ��c"���k6�ze�N؋��Y�Lڔ��q\F��k�������OLc��<���r��1���r��x�{*2?�҈� �Ϧ1��&&+R�FW*d�TxH��+�XdFD �3��$�>��JJ�Z̥��J;�k�u�e��j f�[n'r��MY���[�KQy�A�\R˕�^.�$r�� p���$L��k<��f� ��dzZ%�!�*0���{&�$w�4�e��=_�e<YZ��D^J��(<�rǚCf�n$һ��P�8n�0��I�V��Ř|p[b��L�L5�H��l�]YՀTK|��v����!���<U��H:�ڢ�� �L�ê��TQ��X��3�s�J]`g<����� ["���70J+*��Ǌ����r�
�����8�" �ɓŉ� B�_H���L���!9c�9t�i[H�Jcoy�܍��Ͳ�uo��*Q�;1�1!ś���0g�8�^��VeS�����^\��X�B>S��\�t���V\��2-��B�'�Y�
����U���}��t���ξ��Gv�E�V��Ԏn���]��7�t�Q���I���UZ&��H���X �̩d�C���� ��~��H�rO��� p��3'�7Bv�I�����fc��G�?�5�n�ɓ�mrZ����W�*�;"qǨ:Q����g,�Zl[0�����mZ�v�y�e;?�zvO��d��*��&�cY+3%h��%G<�i`���[�S��ٻ~������^�Y��Cؿuz{�z�b�P���'������Z�.�jj�ׂD��/�|)7'A<�S�꯹t(�He[�D�%�O�խ��}r���+4m�5������+/�Gi�� o4<�V�;�%Y�`��:OA�&��=cս3�?�֗S�5�N�َ��,Z�P|=LfO'�=YM~�T8�7�� ւ��5�jA^��,^��v�?n#�=�#O�G����Զ,'drМ���1��#�x>�{����5^��<Υ׺�;���W)�u=kP�l��X��ceǚ�"p��
'"�c�W�I2�ѓ��[�|�~���?��M<J��0e�8 =��<�뇨�c��W�J�y�JK�@ S��K|����}d�ح�T�dI�zW�o����z���?k�9��G:w{<C�� �&�:�J��E����?�>qV5㿝 �5 ��o���N�BI+G%Y<���q��{I �Ǳ�?�Wi��"a���}s���gJ=���]s�R�ԓ/	��	�dciK�r'�~o
ڇӇ���U%��i����{d
��� a���|{�}}��T�%��{���H?�� ����s��)���Ƚ��ݣ����u�G����!A��^J�A���9m�o��ӧ�s��<�x�<J���&,�%X����*�#�8� ��8�JV��e�4�c��<(�%���	�W�J;|$1�Jyq�e�(�x��_
�r<�k��U�Q�̜Ƞ���uF1�͍�9CΩ����n)*�~ �S%�k#*zcLv�3HG�#.t��ͳ#S�N�U3jC�>L��Vc#�6<����)�XFqVWO�M�g2�fG�s2�K� Ŵ�!��c.7�`���g���H�J�#	���MAv1&��C�>98�	<t<�1.�Wĵb֬�q4#�7�1�e�9ǳE�5O$���� �tT��X����.ɱ��X�<Es)hW(��j<*�����^~��ݒj����1Ѻ��ʴ�����vg迃X�����}�0f11�k+�\[d\ypN,�Kea}���	, d��Gٌ��ʽ�c>Q�(�x�ի�F8�7�L|p:���q "�2Z�:=i2��d��(�fv�+]��*'0�s�����Uq��L�i����J�n,�EV,(�g�;�r~X�S��%Q1��?���{�UŴ����K�� ��x�)ҩx���v�v�����B�)Fmz&�������W�1��E�R�|��iQ$o�ȹ
(᥎�����9
\R����XcŃ�),��8W�nre�l����Ap&��N�p�l�G�)�p�cx%e�*�@��m�Yx��Dded���Uc* �(�p�@yy���f�E��Y�l�w%�6Q�-zc#'i6���U�|��I�V+�m%�KAK��T6���dR�ō����+$���fE�S{�˓��4C=�r��31�h���i�ş�?����2+��d4�V�ZY���e���q������?��K��W���62�B��%��YT1��x��o�� �ʌCL%rq�Iĭ 7��c3P �܊�/��t�篐�5���򱥎C����r�.���,CP��ǝ��i�.K��Q���B�(v�cO��>PAuec$�R
IrAz��*������	֨��~ȧ��#�I�&B�xc��h��r�xl� �!ݹ��:�q�;zc 1�����M<�h։��q�/�^A�U�i���'u,c�敻	�Y��V�*c��؎��~EV�8���3W��(�d��nq���E2��r Lc��.�'����Q���E�!J��j�$Fs�*���Jj
�����Dhf-� "�$%��sh3^�P�e���'i�E����c$�R��&�8�l)�Ek�G�.R��U�QW�`HcHV8�.yj�5˦`�I"��J� T�B��J����p�_�ߞR����c*qߎu���n��F?�b��[.f�ǓAc<T�gP���A�f��b��Ϲ�3"-���$����%mȅh��1f�q�[��YT)R��cp�C6c%�Ց�&��@�|z��MP;=r2ҳجI� m��� b�	q���FaJ\0��c���CO��'JԼ�Ȩ�E�ݘ¤]���k"@Eʂc4m�k޳[Z5��28+P�.⡋
�*��9"�C�ޕ��W�jF�)M��Iۙc��Q�'fc���Q[F�zdc�?�1<|v%)�Zo#W�mʣ�0��9#B�7i��7�*�3-т�΅)e�Fm���v��>n�Z��nIg<L_"6�L�(�*E<��I��,R��cc�j��&:+r�h�d2Vqir�Ɓ��O�UY�Će��2�c"$��:����1;Y@WEz2����o�%�6e�D<�#�&r��D&7uM��W�}���E��F�P&�z��$m2�Uxѡv��˅�R�F�X�0��hT�"��梼�#lG�u���X�X��c	�ƛYc5�C&L��V�i:���y)@���F�+1���G�Z>SE��}����3��j�*  �ӆƋBQ���>qKy%�w�^m)�U�%�C<;�ƪ���sVj�bY��E	e�|�dRТ@4���<�J�AZM�W%v�_�[�c$����4��%x�֛U٧��2j�'��E
���v�c#�0��嗀D�VoɃq�@L-���-\m��m�j1���H�4Zo'��㔕��U+����s_�p'3%g�匔xQ|�_��|�\��J?�B�n9c�)�H�ٕ�@Ō(g� �Z�&ȭCE�h�V�2�֤��vFm�/�2
�<̄0�q�'���-F�W���/6��Go�#�1De�,�F��E�u��T��]�7fT<�X�����0�*��؉
p�����U/'`�ŭ7�c@h�O*(侘�^m>bW���\��58�Ý�[pw*W���錬eczc�"��ǕL�'v.1��y ��~��|�����'*
����6b8�r��֑��@� ����?��N�k�#m���ebN�	i�v <�ln�y�rYH]��?�\d���r�Aqrv4z/�* �0�>��+Ş��o�D�	lhd9ƴ<mX�Jq�LS 6F70� `��C1��J��MiXL4�\�e� b ��0^|�;���c0���	����E��e�Y���䓴؃*;.ʬ�v,�q"�D�����&���(�G4!�]�(hZl��y�cH�c+���)6�2�,��C�jMt*� ���Z�e ��1�HMRH�2���#���Eh�3��+Zj�H���~�0݌���f+�,Ա*�#�E��1�@��s��zc1�c1.��� ���|���7R��F<�!Gi�:�J����1���}����̴�Q��'P���6�_ƞ~�"�/��ʧX�Z2ͱk�/J�����K�hE'
����h�T�Đ� 5�Y����� �JJs�K���%|�͎�*��9+|nޘˬ�1["�%�9��3dTg?�����\�ц<��U8���x��^U�LVJ%��j��P�Vǰ~�7C�JKL���Lpfo���Q�Z坷��$e�������$;�F2<�-��5eȬ_��ކC#��/��C*B����� R*�c劬��ԇ+�k��JdAr1iv\I�F�w���%o�n>��e�2�
M�[`�J� ���@%��+JQ�)�"���c
Զ;^bJ�x��k[�U��E�i��S�ȓ�u��*�MYV>6�[%�1)��ũe´�\$�?���x�f1�7�E+�mT˰y��!���C�\�?؞�c�b���H
�:�|��t�0c�	ɣ�\H��.镳�+��x؅�M� � ��iM��(�q�x֪��!��!����ȼ2�g5�a�,a�;��r�q�:PH�̮\����R�*���ANLc�V	�|ҭa�,#���y]���S�r�����c9+�@�Z;d�D�ދ��=1S,��ITf� ��|1 �1�|KK<�"k��\KI�į�I��oN~A� M��$r'Yv�K,׼j�f��?&*���PC��}�ܯ�2_������Z�G���u�c<U"�!g ���-�)*�Z�-eå�q�rHjU
�s�e0mO942Q���G<ٌ�B����Kd�K��j
�$Sǒ�т�C�:(�Ic!.+�f�[^ƧϏ[!zϓ�v�0�e�P<J���r%X�q��Hc�Q{�b�*V\b2������mD^;�/U⁕�f�ɲ�3$%q]c(檤� ��r���S�*���H$�`�3�d3��Y&B�]��|�����o��<�_��՘��֥'�<G��#J*s��/�@�2`Ы���e'����2y20�\�P���"(��+<e?��E*���0K
f�(�\�4|IJ|�ܳ~*M�#2͋;dcTR0��8)��e>K�,gnM���y"]Iݞc�������P��6��ә!�Ҥv\ �R���I$�%��c�x��=�W8��Uȥ���V�;�?�Qk�bY��f0�r��\g��qR�+8�^t5�x��.�y��i�@��"X�.w��RS�X�,����h�iV����1�9�� OLc�z3S����0r�3ꭾ,��5w0��\��M�n�J(GPU�ٌ�����wh�jhSm��Ʈ!���53�Ѻ��3\�1�5�3�yB���	��K��j��pU�>�.@T��=�~=rr��@G=�d~@$���{�{����۷z:�\�G}�4�3��6WOjխ�t}5}GM{d���Q���;\���a.���F!wg�oUˣ]@ִ�\
��7b�eBYWrJ�ǐ*���we��0j
�ˑ�k����Z&T�E�yq�#�rg�O�.��w��;�����7=k��#HЗ/���^l<����åu��E��?Q�ѱgͮR�<Z#��7I�"ʑbH�����;�n [��RO��M�S�YE(YZN;�q�{��U�����>�����K/������ O=���->����V��0ݧ��w�VP��}Yd�ˁ��p�J���So��꺣$��
7pD$Ep�ڿv'�.� Q�@�
hi��
v����ۏ���U�	9��Z�4�m�%M�T�6�Y����޾+(��9���>��� �zK!��_c�<�l�#T���_�-�c��@��RsPP}~�}��������v�$�3�����'������;���O���>�������03���)�B��0�?����e�Fz������(+�ۑ���Ҿ��ON�RĒMBKG�#.�v����s�?��v�h|b�DTr����G�����c���p�����GS֫zQD5i�u��aͫ$�d�-��o�V�}e�Oԥ��EVJ�Pp��1<��n;�����VMɨR��IgI�c�U~�������� 뛅�Y�N���y�p��ח2ݾ����>wԹ�u=SUӛ�6��	oGW����x:K�m��=/p>�j�vJ�>VH�Rf�b�+��Db0@G�f<�%��]���;E��JV�nud{��8�k�^�i< ��J���{G9���?r�G���۷���N����t�=_}Aum21��Ez�T�5�'�,�/�5��Z����dg|#톎���oK5,y�[6��|.k��%��~ػ�`;r1N��\�[�f�Z�P��F��[�)b�$O�R�)!B)��e�����w��15��zL:�O����$�O&8�/�t��bj���8e<�B�	���6����M�+�z-��>��S�f���@��t̓D���x�9���'ďN�<�����>7H�`�v��h�K���G<(��@$�	����T\MQ5�5�l0-Y�\G:ľ)�ӌ�V
�˅O0V���v���ɽ6�|���_����N>�eQ����>=�E�6�;��/��	c��_�CfN(�nx+q�Tv�W�c~}G$ّ�%3uj+�E	\k������Y�9�G��|�X~�Ǳ��� /�mW����\U��>*+����Oĕ�[F��(�-� �Z���~�1�8qe��qRc��b�hd����@.�%�gSĿ%V0ɒC+䱕f�s|:^�˟�bɌ�<x�?n�fQ[c^%�'�)&t�JVEp���\P1���*�"��ȓ��`�a�1/&pܗi�tD�7��aR9
I�n~���y\���+������c�ex�r�jOzb�n
��C_ΔlUrg�WK���r�"�ˋ_ ����fz�����G�7�ఃc>+I���?4�rg��C;�n.�(J��X���u*���l���K���b�J*�3��H�j1�5���C���e�(wW6��ⴔ����r����1<^[��VLx�KD��"���@���<dKn\G%#p���b�[��g��$[{AZ\"��1�Y|��Ԡ]�Ef21ÛJ���q�|�X?�32�ǙΜ�lG)�_���c�%1��iM�Ĕ�]�:M�i;�U�s%x�@@^N���1a�����2)�\�ǅQ���"�l�VE4�D���R!��F�C�U����so0��!�|�
�n�ޘ�A��JfZM^4�c�����cLJn���(�%_��0�W���x��,�Kگ[HЅ�M�<�h�,�X��?ӋL����a�Q�F�NW���[��U3P��5c"�Q����uw7�,q�#�5*c�ٕ����@��;!QJ�#X�g�A��\|�pe����R��{���f񱟍ˊ�1�2c:͔Y@��9�"j?�:K"��A$9P�� 4$�c��=\�=�)b��joQ����b�S���X��Lx�Y������,9�r)t�@���;'�(��H�wb���&F9���O�ƙ4��ޛ#�2��
)I]��W�W,T��|@�*%M�!(.q�_��F�p��`�����e�
Z��π���d�zb�ǒ#r�����-�c"x�2���|zy���9)e�,9R J�6 م9x�2B����ѩ
W�d�� CzS-ŠC]<�]�+�/��26!s�53����-pם����&�96]g8���!�P[�x�1��Y�gd�I��d��U�Ϟŕ��	��Y��,`�XW#���|�U�����2!Uj��A���|!%�X�����
U����zJv�ٮ��Ê��˴�Y1c$j�N�tWV�b��)h�)�g�sV
���"�!r�����䴼�:d':&4����゙��o��d�"g?;��\7�L����$�c�����(���E
k��P���F@B��+Ù���%�,�]��?��TP�b')�C)��'/>E#���Enq?kx��'�>۳�0/�t��NX�r�U|�k�/�N;�L���y;?d^}1���qcaj��r)�'�ȿ����rP *� ̵R�$vd�~�	����9c��]"�9��
�+�eb+��37&'�K�s�6i���$z�gdV�(d4uBK#m5��S�VmLWn�����I�
W�-J�B��H���c#�\����/,���&x�x�m9�E-!�}��>���()62��f��q�1�-|����¯'n�Q��CAF�±�.��s�.ròw\fy��P�3�-��(�I�b�C��Lb.,0NCf��t�:_77���O���?�&���%���L`�d@ɽ��\rM%vh�q��dx��5V�8Pqtc�k���3��*R\y��鲴W�3�(�Q��P��Ac���Z��_ڄ�k�K<�^<�j����jnɻ��c���PU��*��1�ޔ�^�b�ᤈYW�\,٨���2�%[d�C5�M]���MSN��ȧ0�X�#���
�'��Xʴ��E�OX�j<h2
�]�H\�����S#İߋ+���� q"�Բa�)�UXq�+M?{xPL�F'���bdC�i%�o�y��3���<k��ĭ9���!�;'�2FmY�g�
l���T� �c�sS:
ۉ.�e�Q �<�d,�E���b�?D�X� +e���y#DER6!��w�c�N�d�<Ҵ�	X2�O��.얝�.����+Z2�ظ43F�B��rXy_���4�P���Gfa?�_�����i��$+�YR�ǈ��Be����X��ڜ���nL�1�c.V�5������5���to ǣ�7�K�^V�Q}1���+{��_��9$!Pi�=��.��X�3Zn��,c���i-_�L��x�rz��-����͉ob7eUe��$kI�i��\�:7'���;́9\��G���c(��U�3SfRvm=���sgyq!j�~5$�;�
�7!q�<�c�'�|���*98Ʉ���ɃK~M�$�f�+ʋS�L2�=)A�gۇ�P&�Ȋ�dM�����݁	1D�I�^��#�(�ŪU&%vS=�!���1�~�I��?�j��Gi��D.�Z����wV(ܨ�[�t�����S�IV�fȫ7�򒁎A�nL��Gezc�.>��2B�(!x&2;m��T�ab��-���W,c�'jھ x���7<,���f4bq�$�QCNO��区��Q
j�E*�R��t�)e�����,>	��Lf�US�=|���"ؓ�Iʃ��hE�Lq�ncr���̖��>������i������u�!d㿑[��.�q�N���2L�'���D��7!Q��
�Z�%����DU���аc�/�mx?�M1e��DKd�E ��E-?���)��2��q_���j�P��"�E�g1�g��=�[��uU��:�Q錍�6U��2f)L��_hɱU!H�%��guR���0P�O>0�Cc���f�)��(�,��sVF<�ُې��e�F7t��δ8�L��N�isH��%nD�<��9�g��L�T��M���,����90�� [$�.9�y|:m�)T
@m�1�CHL�)�4�O��lcFQ�2��8�9)K�[?��c����,�-�v��'�*��1����FvY���!�!�.3DٞU��7Id%��%Z]g�9���!w	Ò�m�1�6�J�vg��+��?!��PO�,x�j�X�;�}1��jr-����[��?)�J�\dYQ+ �EYxq؁�1�c+L�)Y��C`:;S�q(~d)�4����L��(FS�����3�R��<sS%���I�n�;b�����b٩
�(��Q�,2CWP߸y�R>˝J䪼�N65��ljڦ%#"e>
�d��9n
���2Ǫ6m�';#���&�p��x+"�tE������0�<\<m�k���d��h�+6S;,�eR>Z/(J}|h	�b�&4�l��iG2�⵹���<�)q�W���ۃ����2[���s-HZt�R#(�'�Y+ ,'���8�)��Dʊe�W�H�����-j������/2X���>�κ%!��Ǫ���$ ӚV~<Z�<� �,G8�1��«�2��٧I�T�F�n�raH�a���Q��bG������Y�.jI�cX2�Aq̭v���3G+0��,�CV���ě�i���M՝r2r��V��9� P���r	\A��㡤�t�4%A��V*��ڒ���If`�*I&���LeR�0`#!�2 2�+��T1����C�=1�ah�Nh���kY��-j��52Cѝ&��%�#0�gɌ�����)��j�O%3[zE�D��2���0��Y�zc�� )isdzЦG�13��'��yl���1�ŷb������a���aX6ՆK��j�jHE��'�!��T�X�:l��1�+��G|�?�^f~5f��U��Q����Q��ٽ1�=r/It�zǺ�M��#�IDF��5�M�~����'�u7�MII�˘�,��޵i�ʰW��#q�Ó�,~ʿ�>��I$2H�~O���O�g1���C��S;Y�{ql�G�:oHԲ� �N}�ԩ��R�?��d;�>�h�18>�RLV�;.@����[��W����bb;H��*~�f���H6)5��G��EAH'��~�ړ�_����X��}��uݫ�.��������4�;F�<yiF538`u&�J���VL�3���Lg����܏V��n-
�����9n�>2���C/!��U��^A%��ʪA�[��,_�2�8��>�o�9ҝA��d�|�
=[Ӟ�{˛��R�:�S����)�y����}XJ����S)�R�%���l-XcM�a�-t�ZR;��9珥>��8�>;����]%�Ks�������r� n	p��y��c�:èzߩ-��[�Z�W�^�ᶡ�kyg'5e4o��M�.&��\|X$qq�c�S���D{�t?~KIbx�O��߲S����! �8ǯ_��� �9d���j�k��5U���@�1�y726�!G����H;l�#��G����o^[2�e�}�?O�˧N>n�%c���V9v�O'a���w�O�&܏_c[����U��e#���#�~3�"`��J�}�}<��-s7\���&�ش��V��U�������f�x��܍���,([u�?ynI�7~���N^Z�*��~2�x �������7�zN��ί���VJ�¬�kL��̎E�E5_��Z~�<�A$z���oO��V���qS�}�I"����~�<\x'��oiچ�byt�XϮ��� �>���=� �5~�u�^OH��Ai�����t�kC���+�̧��
��8���Ɣ;���=�����ƍ�%�c�̏�dv�	X���~�`s�V�_UӦ��4Q~��2�(����z���?L�o�U�]7�_r��~��t�.���kz��x����a���^�Ԣ�9g��Ʊa\\��J�f����� I��KoհoG���z�j�2�B�6�Ơ��W���%�H �:��ɶ�n�t[U�7+ǤՇ_z�& W�Ph*
`���J ���B@^��7w;��k�����ӆ%j��VQ�UZ��*�������/͸5f6��vh�k�?i-�+p��݅��d�@��>> ����Cu�Q����.r�9bXш?چ)[�<��	~�*Ǒ�C�m۔�qz���,~ޞ���X���#�^��և�O��]+���s���X3SM|6�kYFC0t�毼����:�[�`���GD��)�{�'$&$m�+`?�����{~h�6F�����J�&�8�FBڣK�׊���s9����<��[8�$*�Ŝ"+p؂ꪴd��^_#��� �z�j��$��~��9�+��v}*O���|�9�}�L;'�{�뎖�:���;���z�4/�/q��@�z�8�rkD�:Sg�5qr1h
m�'i�<����=z� ¶��_�}ֻg~F���(ؿ�}4z�z�����F�H�[1��χ:6�JX��nm�"+�WY�)D,9WӬ���62y"��)��ȝ��os�1��.��.���w�����DKH��99�?�G"�zƝ,�	S"f�!*���zѝSn١Y�JVa׶��2�T����jvGp�n8e>����n���N�������i�{�#�cw��11�{X�ѓ��cǴ1Mi����Z������s��"�į�����f�2�Q�&�u,�Q��o5���UWh�Q�T_�T2�S�>���<�jk\L�ŕfŹ~ä��I���p	��~�͌��<�*A�Kl�~al�_�LYa�[���@K���ш)錅B��΅f�e�!1qȥc���O�����Ȑ��S�6%o�t�Ӊ�G�sqQSu��y%4w�YJT�[q�U������S���[%�NeR���$	�^)Q�fHRd�䮴F�zc��&t}2�Ѫ��#!��!�F:��AUT���4��&3��k����9��R��(ҏ��_�cG�R�,Y��S�sU(�V�2p��)��d�|����������!%QXɴ�B�8��h��>)y�ܣ�(2������c%f-p���L�^[ȹf� u��zc�~5�[n a�?��28f|th�R�o<�.D�eLv�t�����#Pb�D�:����q��N�-�V�E��I�ȕf���"��*�6�� ����ZOl{Y-<U��(���F�����EV�c\F�I�?��i�́�֮��	���&����	�8�g��L�$�aW�3c!JҴw��ʊ��*�̬eB��vlS�Z(�˦l�����z�T<�>�Uأq྘ǳ:S(W!Z��ѲU"�ʅ�i,B���l�\'Շ����j�x(>���X�-;cB
�4+Lz��x�����o���}1�Uʕ%�P�P��X�. hQ��cB�P`��K�o���Q��t��'*~T���	�����ro���R����vc�J�kU�qzEL���B���JeѤq���|3	���x����Ή\tAO�$��E�+JSM�4�7��e_"�匵ZQ��ɮK<��4�ű
�O"Vg+�YG���A�&��f2瘡�?n��ΔR8	ڛͧ�J�ii 4� ��hHV1�W���*�A��y��X�=gz�Qh��&�n��Xȕ��Y`�Q*ݲ�ł*ř�p��Y.E|<��*�S�b��X��b���v�2��2�(��9�E��M\qv�GĬ=1�(�-���
1iX��J3�ZQ��)��3�j�P�wPX�T�n����=��s�&�1O&�Q��� T�9��:�t��g��(���E�,ut-h�㪔f� ���M�1
��,2n�GHU
��$�'9�)<x䤦�V��M��R�}y2;~=+���V5����~:��N�ۆ�R�[8,�i�C�'Rյ��
kz��Z-/ڕmDِ��u尬���b�,��F92��`rrO�%i�4H[)���U���Y@^ALa
Rj �Er	�Z��y��Y�f�h��3;P�>��R��	ƙ�ęd�{����unc��x�+�� G@cl@�u��Vr'R���@�0Pȵ�?�'�m��c-��ع�DnQ���<�R�O �T��K!�a	W�E�7���ӅB���)���mf.���9UU�J��9,`*���o'$Y]��	�7�'d���Tz�Q����6����2�q�'Z�^�s8�Q9�fǛl(���2'fb%q�7�"�@|2I�,ZѲyq��U���՘>ĄR7R��3d��-x�[&L��%��j���l�x����@P;2�c*�����	� ���*�Z}Xd�$�W�	��Ԯ�eA"�*�Pl���+�W��yܪ:Qf�`�ːev0�Ⅸ�y`O2)X�%G��! ��(D6\SA��K�(%���7`���1Ua��ƌS܇>c�d(U��)6W��ʪ�/����b��=׍_����Y_��dE񷘃��;N�B��d�����LegM�q��i(b��p��k.N\JX
�)lte���'�r)�\ ��x;1���d��j@��o9�q�	'�Mɡ�� Ы9�Ǆ�c��æ����V�&r��b�wi�qϋ1�Lb'�LR�*�9n�9�dޅ[�d�"�T%���˟�;1�'8�2(?zq�:TEҵPeZy@L���B�P$���]Ռ��-iX��$4�1Ғ�W�<S�$�U�������1����s�2o��q|���b��C?�@d}1�~���R��ՠQ�D��_Fw�g'��p��1V��2[����Pc��g�(Ͱ
�;?��*�,d{픥җ{�{RW]��'	o�-~�ԁ�p�2EFLǝg�����G������VZ��\; ~�݌yh�߹�y�����#J~�mT;-+0�����;l��OLcM�଑�<1�D�o䧎�Y�g�|ՙY��g���e*-mGy)Eǚ^����uE�m�2�+�d'��yw����#5��"7�a6"�' %'���e���c؊Y%)�8��1l�E�V1�1�\3�%�!�>�Ŭ���#i�qiW�V�PY'�b]���2���>����Dln1s�b�#KZ�%�cHф�Ra\)�M��U���HM2�'�<�jy6�7���AUZq*�-�2zc&a��(�ĩ�K	�L��1��ʥX�*)�U�VM��T1�V�эt�%�6k�� &.��?;|�Ǧ3Fs�Cc�M�N���qj�!<0J�(OW����,ĳ1��>�r���<�6��&�&`M22 �t+�yD�`��ĥ��M�Š�ԡhcy2��e�2�0g�Rg��oSU���v-��#&�-*c��l�suq,�o(Vx,�2�,����oLar&�s*��ӕ���Ru<�&�[lw�z�H-���c*��3T��f�1�d�U�[�#�<�G�p�ه=��%�������g�R�3ѽ�=�� @࿸�<g��?���lŌ�|�7-֩�%��[r�]��W�?�nwVn[v2�e�)����]�J��L��0��T�[�T���§�~/�kW���abؓ�G%���1��0T��J���r���Rz�lwǦ*R�9d
B,�K�><�2 -�p�K%�qm��	3ͤ����&h�]3f�F(�B�r;(R�d|�N!0g��Y[)1�9��Z�Lg;��ѣ��]l�����8񤸌�N+�eHe�O`���#�*��AR�غ8�M�1��gK�4ɺKN��L|Lj
;Z����%�|=�L�E'��9��!EY��Ү*���j`]KX*�wfLe�g/*%�L͕��IyZ���O3��)VdVS͸<X�-�*1޴Zp�țKɃja�szE�W%~r����T�/��#��m<z�IP!$e���d�HK�yMb$?y�"HU��M<L��,�Y�����%�d���;�K�)0��T��K�c	�+K9�ƿ��V��v�
�@����rv�X�~'(���ke�R!:�q*p��!a�����g�r���*��8��0�4���Z{�7���i��`��y͌J"A��K-\N��_��?��O�aC�/"hV݅�1�1>X�;��Ŷ2#���N)����_���X�c��Ԣ��˚�3�6N�F\�����՘ �����C�!�&�����ў3�_N�ɒ_�#���(ÐR��:���R�u�-N �1J)ࡴ��=��UU��R��m���26�{fV(�h1k�3eRA��)��^,�Vb~��!�4dd�~y_������զ3r['��ג�?<e0	�X��C3	%������+: ��SY�g5R��±�:)m�yg-X�ɨy��,�g�7�3T������2�h�����	cdd��E�6"6F<����� x|p|�	a����c>��j�i��V�\��'K��tm
��t���r�	��/Gw^��C�L`������7�q�d^�b�Y�CZGE�9��`��H���� ���ۺ�uC*��#�
��IIW���c�3uw���w[�:�������7�z�X�:_�:� �f���užFU��N���tl׉�)��qERi)��i����@ø�ݠD煔8=� -/�9`�))�R$�i�'�<��ϑ$��G�.�Z4�s���=�����Yw;��N�ٷƦ�ӝ���+O�����Nx�+�='��4�_��c��X���.u��ig;�U���ݟ�?�k(�����7>.Ė.	 ��笫J!H9b�0��Y�H^o<�A�5��~�5���rz�p��M�D�Q莝�|�[�����.�ub�Y]�ָ��H�m����3�oZ�5R�;	�{vF�zT�ynY���\���V��5^�#��c�� �� /�<~3Z��T������27��lC;���ؾ������E�U�O?c�����T4�Հ<��?����t޻���3N�#�26*כe.B�S��c� �5m���R�1�8���/�r={<s�-N�@<��,�������?��=����K8������җ�VC�6JN�V[��R�O��l=Z.��NXTk;J�w�_��׼�� X�~`B�D���?��=?Nhw�!�c�ds&rT�>9�Z(�ERh���N��'o�U:rM�lIV�.	f�C/܁�߁� ��.�FN�=���s��x� ��x�%�їCu��ll||>���m��M��UuW�|`LUWz4�3[*v��յ�
��5�����x-��e��{��-��r=�1cJ��'�I�X��*�=�_׏�����ꎠ�Θ�����gKj���~>wUc��5G�]R�֭�f)�}��(!��	k�=����ִ�:Rbx�6/<���݇���A��J�u*v4xa��X�]�@�4����ހ���{���]7�[�=����s��j�M����:�x�����4Ѻ�W8���o���zn��j��e��0ƭ6��ѳk�rm%�y�pjZ棭�_Խ�R���h���<�U�	�d���A՛�<fԭ��,:t�ZwM�#�Fi�w�*#��R�������#�;���=��i��=�����~�{�B���ǫ�񺯷=�ԴD�������u�k3a��6���,{�y=?�3�u�3dj��mֆ�[jl�n��;S��P��JM��e�M"����?x'�E����� T��f��8}�F�H��ݮ�N�H�F�!�LKz���?���e[P�C�v�N�!�ek���.��z�Xv��/e]��/�z�"�h�����8=��a��(b�p�mv�7�L����~3��='p�22�w���G5i;��uzȆz��പ$����J}y ����g��}@նv��y6��b�c�Xh���V���	�H�^S�B�/������]K�:oC�#���ӭ|n�к��������ꌾ�ȌzSw����
�DH�Y���yt��.��]KM�6}�ߖ��E��	E�D-bV
~���pKv���vT�����'�5-gx��,�q�3����-���O�Y?�Π��7�U9�/up;uێ�n��H�]o�:7��U�O���qu��S�&f�������r�<%BB�UŧC�b��Gr]���55�b��C�DN�N��g`�ʏy)��=�^ނ������Lv~N1�4�'Y;.�-�~Ҭ��f�K*w3k=���ڧ�=oC���k��z���������\u>@�]-<�jX���9��G�s��*�&�ś���qS��W���=O{IE��h��4f����D1,b8ު��"(� i�d���؋RG�Χ��@��mKpi�n�%�����e�+<3�R�,$%|5�r! �J��z�� лA����oRu�o��i4�\{��n�~�mSP�4s��vζ3���WOǽ�mʸ�J<��}!ٚ?�N�յ.�j����tࠚ"�Z����=�Z��C',��4��3��v����|�?[�L�z�~Ϗj_�U�\o6�Z���
�
�� o�ČObE�,Q>_Q�7=�h�F���]����;��Hd���~��������%���k��5ר�����ʵ��s�}k�����5KM�{�6U�/kտ-K�RI#�U6*Y�֖�:"y��� �5�l����u� diuS�Ti�J+n�Z����8n!�R�MI�RX$�� J�.h>&���VȾj�da^�;"vL�;c���3��χ��X	�r���b�f��{�f�?��>�>�x��Y���?ĵ�R�X��e�� �9�m�۶���5m��ì���&=�����.j�)�4S�8 ��[FrU[ytl�5#k�=q���*_���ԅ�ǳ#�P�m�A���b�j�v��L��\��Z�z�0�<*Քm���9�=I��e���o�$j:�i�T�c�a����rr�d�FTUWJ� y�s���  >���~O�`�>�}�����?9��4��7lc�[-|�i� �U��q�!���D4N��V�P6�錇+�̸꘾e"*&��XL��Ơ�9Gfc2ȤtZOb�*�2U��L��[ݘ���6sOy�q%`�4<²6�c�ZR��O��ƴ#*��6UI���M	�UݶT�}1�i���o�O������g:���O�q/gf-5�집cLuĹ�%���b���h��h��������D����B+1��88��IM�V7�yc�ފ'%y�H�&�WF,ԗٙ
���Ǟ.��ɑH��e��,��J!8���^���1 ��\�^�T�c>k�[Ά��䬲�Q�X/b�Es��8���YF#W�6utL�wb�2��j��t����B��4�3��*��:���K����bb=1�W���qi�����*�I�E�BA.h|����̌�Hc6ǭq�d��'��鵖���&<��Z�Wr�E��>0�i��Q�� jn��H�R���9�5q�ƃ�nP$R#�@~Ic$�+�mZ��y�6Gʂ�<�
�vi�,�0���c���P�;=���|����ګ�ԚR~@X��f
���W,�ߏ��vV�L���	O&����)�rd>� �����9=��
�ȥ"�Ή5&L���`��e-�E�b�6S�ˏ����%)U\�Ӏ+����BɹNswr����J�]�ES-�jZg''#�)2��z��Ƭd�<ʕ,a�f9i�U�1�9O��T��\�.�m�g���er�F0P�ō�fMq�!9��wy�ДkB�� ^K���wfP*X�s,�����o���)���x��y���'!�d%AU$1ԝV|�##�g�2��?@�|��쪣}�ҖR�0�<g�%.��[��ҫ[46���9�l�0�=<�J����3P���MU��d�cMR��Z���]_uY�+r�����]�ú�QI
+�J��F-�I�҉ ��gu.X��zc"�o�FTsq��!���|��T
X�Ѫ�IR���cE&q�  �ƹ,������˂����MC� s
�La�d��,���<�	���vYc6:Kb�,Q�bT̐���UNޘ�ƦE	��`�Z�U��k3
�GlM�4f	902��6�K;,ύvǣ�2�)'�3��<Ч� 	9T!=1�eI$��>k�&�&�.DZKt���q��1�T(g�0v�|�A�z`Z����8�<�
0F�ܿ��J"����\�1��#�Ԧ�-�ZIDl����"lF�X����N�|{�亟ɾ2��R�$Q��ɐGaD�\����_�R�c�Ld�>NKYǐظܩ�4>)b��Y4a^����<i2�g�о@8�<����`~&�o�v!#fm�Vc)�f�LPUnJ���4��B��kS�3�%y�`V�X�Q�l�eg��c'ǚ�O<G�����d2T��Rʔc)����{�!�K�gM�̚��b��A]��b6�l�*�γ���9~p�2Z	�k5�V�c�#�X.����
X��wE\������D;<ryB�� ��� �m���<[ c����>4��	%�+J��>%^%I �6���b�I��6b6KMV��cGi�x1�'�(#�ܱ����K���KR����.�U9M�m���Q�C3��3e�\i��re��$��5O<.� �*��ܔ�!��(��'«7|��l������iҀ��Ӧ�YWj�%�)͌ySz-�\��X��v#"F^O>Fɴ�5���&��s!���Eg��N%�%�����jQ��&d�^L�q�`��gA�#����,��9�ƀ�hU�K:�q[���0��=�hx�"��*����2�!|�9c�v�B��l�;���L��@����#��C�^_�[$٘��Ո3�����f�������#��:��`(�늙AU_��S�W��͕Sb��M@>��<�cp��L�Zk2UZ+D����
L��p(�V$l�8J��j��y2�[")�3����L�:/"A�݂�5�D�U�he4�R��|���� s~�d��I'NG��p,�!9~|ޯEy�ӕ,2^h�j9P��Bm�2l�l�R0�R�C�5+zdʈӠ�m�^���q�|�������d.<��"1Ƣ�����@�\1 ���$`W򦌗��aUgc�3�WcI����c�y�W83)㷦1�ԋ��#�c���33���+���f���Aı�FYQ�C��/�� q|��;O��.g?"����ے����4�qnh՟{^��Dc�}�h��Fŏ5wA�n�C�¿��yV>" ���߈�u���? t]�x�Q��1��+��f��2��3F�Yyvd�JL�������Uي�cJd5(Y,X�(4 ��$�?���������c1tk��D��D��]���?8�����&nej(�,�2q nLa�Zŷ�'�� o>�J�D)\!��� �1nd7,d� ���12X�cJr)���a�
��nI�~A�$�8�0cX�+�Z��c�L�|�P|C�7�^l��e���ʲ�f2fJ��RJϔ]�g�5�o+���9�!eR���	ćc��vZ�eW��č�[��V1ȑ�Q�@�J	�wp��Nȅ*#hI'2C.�D��R�|��9����AT���e
�J\�̆+��ዋLLKc>B��*��L����6���y
S)�߉
�D_al���y�`�� 6<*%�� �D�bWv1�y�rrk(Z���t]�%{))�4����3��z
��W+!O�b�a����7�9�;�Ǔyb���DVc
ؔ���Ew��(%�<o4��0�d�My�0�{�\�����	8 h��6
�p�g%��F�(U��k(sGx�c�H�c®�+U��6�[�Y6@���b�������Z�Y4�fm�yޙo��7ٿl34�h�������_+j���I���Zb�P��K%jI�c�`UYU�˕�eF4ܛyq�	v�՚6�g,@o  (�N�d�mlzc�SK&�4���2�����c�.��:'�*�PA�9pZl`���m3h�C�G"jR�\����H�	��R&a6�W�WU�y]wȬ���9�L�|z"���Fs��wB�6c#I^�	DC ��qّ���1�����	g� ��agƏ�ZcP�V�ȁ6p%�h�X�[�8�"�o'��0�3��:ՃA�h�4,j�$�ygQ��$�~E�VL��X��?'�Q�,��[e]Z��Z�2�3�y"�x"��w�  1��Y9A�I�MR�v��C����&�]�{��+	�X�j�X�a!�K��gDeD9!��@���9II?���tb�zE�q�Lm|э=�� ����Z.'�Д�����c��Ό�I.M1ű�k�e�#ݩ��h� ڄ2�gY��1��3y[��'ό�*8�mZ$!���$4e�?(�j���c_�I��.�[�s�K��EF��,�!4�z��Jr��91BqI|��3����^Eǌ�Lŧ/���~�����V����n:s�m����n��d6̦0����D���T���R)ř�I&Y�e��V�ܾ��$�� ~���ω$X�����s������д���:���#���Fh=G�F3�l�;�tά˔׫ i�:�аmls��5_ü˨���Ƕ�
�bv�f���{�(e�U�Yy7R៴�2�9�M�:��v�[��?I��-�{ӸU�!�� b�������;[�[�5�߯2q��u��^��[P�A��6��e�0�-{E��yI�ھE��_���Zu���*{ȍ� �E9��g���B���T�}+U���v�VUܡ�}�$����C*xn�P��Yh^ܺ_'L�:�ܟx�5������S�'o3�ucl�^�h]C�r��ԟյ���Z죤5��ҳ&W�d�lMU(G7���p�J��>�^����^�sٴ���ɐw �c��>��`��Ï�q��c��}O�y�Y�:�Xu/S�}]՚�??W�z�&��w�X)��/Nuń�c0���Ex��x3�cUNO��o_�~��}��w+�6=�G(����� L��Q�r�\	�d���K�I'w@@,�X"*�	?��*���-�'��_��� �����,RZ�xT��G���NE�����|��..�+Q���=uV������� ��y ���"��r������� _Y��$,Ԫ���?����RƦA�q��y�ycm[�0|#�Lr1ʛPO�c�l,¥��O���{�w���??nG�+�LC#�b��~8�3��Gg�����i�4\LH�R� �9>E�AǛ�Q��[i�9ox��}*���n:!�#���~�'�9���l^��:�d��h$����rGMu$�mk�g�t��t8�o4|�PŴ�ev�G��SkHu�h4{q^�q�]{�?Wi�V#���<g֜N�~)�*�Z��n��s�~}��a��Ω׺~FOz4MWA���y���M��jY�h̎NF��Ҹϙ�|@b�I � �XZe��J�u��;<�j�C�!���p���q��rs-��k#Ym�4���J�'pnПq� ��{9�}�����_q����[؍g�;Ӻ��t�d5�lG����K�4���:_���K�7|N�8c�j�ӵ=!p���#��gi�C��[@��M�OF�l/� b����u��E�X`��<G���ⅸK���О������I�֥B�� ��]�Pٟ�$��/k%�t�X�R�U�� �on_��D���uwx�;��a������p�֓��s�.�||Q�j�޺�]:gܿMc�`b+�H�GX�ba�� N���Eϭ�O�n����ܺF�M�r	����c�h)c�Wqi��7��3��Z�$�<�++�X��,�?j�:�MK��m���5�,B�-z�k2^Y�[��'�Љ+MVS_R��'�9f�� Ӌ��}������~�]m���E�L~���Ӛ?y�֚�mOO�7x1z��t>�t����feP�RǄrB��b�W}e�]��Tn=١��Я)�,ϨAb��"��Y��9�:�4��s��n�t�p��7nVE֣�F�i�6j�{�Cm�U䙣Fٛ��� �G������wNv�;���պ�;��ް��� k݉���	�`gv�G�1��?Y�ݨ5���e�5p%�����/\t�?km���˨hOkү�]����oWe����f̱�ҫ?!��k� �/kIODoj۳\���hn]߸.Kr�������p�f�"�mN�2|�H��Ix��,���]O��WS{����N����N�4<�x=��M/��ޜ��]'VӰu-;�1Ѳ���\|g�M:'N��Er��읇�e��3b�#q���6$<:\��%�K�4�K�*4�*p�VYQ4��$M*�#틸7� ��U�u��*o+z�N;:�\Z�-P�ik�4+�������8��-U%4g�{��od���;����{��#R^����݄��fv�E�3+L^�Ɦ{��j�o��Ȥr� us�����]���Mr�]+L�Yf�K<@9!���=�e�>(G�pd�v�U�O����	�Nk�+ D�ϙ��k�� .�<��x�#���WV�1����:������u�u��+��S|�S_�N���֡=SK�k�X�<�%�j���c`�]���6�;Ѻ�&à��86�5���b�Z1X��k_�O`��1��x� �ݗ��!�~���ۚ���(����͍L҂�����$kA$X�q�x�v�ey�pe��������Y���N�����a��B�����8��i��i���mE�Y��a%W�1���8�WO��l�{[`��t�ʹw��K�5�v(Kb;���h��'�QdFW�؃���'����~�3j��H�s��n�,�*+-���XeO�-�HikI 0�'��5{"H���w��h��z�X���_t��=�u�����w��z_�zG3�� ���}*+[�|�i�<5U�A���a�jz��Y�ۇekw���5ji�[֢v���N%�BxR%a]�4�2����&��IV���v���;6��@�mV��kVkc��f��lJA�NZ8cNīL���� �Ok�=����u�G��w��XL�C�o3��z[\끛����S$J	v|�$�1j����������t�DV��׶-=j��*��U�4RƱB	�5kO6����,��1B�"*��tk�{�\��*��փ�u3-�1i��x�/u�\ٳZ�'s�$�(���W�o۾��s�}C�u�H�c����{v˽�|M+\����C�4jd��.}��rR���������Nq>��bꎝ�k�'I.��
\��Y�)n�JP̶�]U���Tq�%k�@S�){��Ӹw�,��h=We�.�;ҋU�^H��芆�v�|�4�2��I>���¹�F��=�������q�����z/Q�u>��r�Æfa����^&�C���I�T,a����[�}`��]��#�^���?l�T�$!��x��^O�H�s��{�D�O���u�U>_t�Xt�'Kt�v흥�_Ku��D���^�wH�ɣ�\��aG���Tռ��-�kG�}K E���Ѱ� ����}��v9��%���(o�� R��G��v��X}}>��݌�Bu���j}m�J�#�4�F����,-/�u�cv�L,=+M�w���`����l��fiQ�Z}f��U����d=ʈ�*����Ï�o��TOD�і�B��
[�2?GԼ��������{q�	�{��~��7H�ƣҽ1��Mk�thjm���ei�n��d�j�����������&ߏ.3l�ը��Wb��Է�����s�]�Ù � � s��� ��g�/�͜�R���2	����f��)� r�dΐa�y�X���`�&gJ��
��~5+j�X��"�8)ه�rX�,�S�X�[?�!�?#O,��M�7<y���Ƀ�Y�aN,`��SdW�V�D�*��Op��� +ʰi�)�RUU�3i*���4�h��("���g��a@��.;İC�[]��5����$Ťl��WQJX:UyD��%	1�7��s�+��1�1j�*�!Q�iF��(R�F�dq��4��Hb�ȈW�ܛLI�-B�ViU;��۷�1��_C�D�ѩmgdwU�rť�XH���C|є'0�c͎F\��x�J���nǍtՔ���we�T*�Q�1��w)���BƏ$��*JY�1�њSN4<6T,��OLcg��EA���/�R?E�X�|��z�v�\�`F�)ql�Z���AZ���(��x�Wc�`�;
1���ے�û�I���c8�G-��8��R�®��1M��y��'�Qh��4�Ȼ��8R�H�d�q��0J�W�=�q�Z(
��e<��j)��KZ;�1ٌ��oMB��&��ǒ-�!~/(�|bl�,��Fz��ȫ�Y�]�Lg#-���f�'-�(���H���I�R"kK5|�_
N|(q�E��)�5!��]�'�2�0���q��J��e5oB���|4�Q̋��,a�f�uQ9G6�=.�E�<5*�f��}v��:��a����>>��p�2%V���<.�rg7.�	}���0L2�+#�gE$pY��'���R����`�2)��Ӯ4���qf�=�7{63"�^�%2�:�
��X�ԶMf�ܞp��hm\:�^oi��3�9`��8�sN<Ic#�*�GJ�g ���� ��\��`m؏�P1���K�8̤���*U�k<�7NDN�<�e�C/��	d ���B<D[!���eV��_7��'H� X(N&cg�T��*�V$
3�#��N4ZN|)�)d ��d�Ki4VTV�Zѩ)\�L��^@���Dn"��@���6P�� ���(ʳ��5DiV��t���-V� �@
 vA�0�e�NU�	,&'Sd��0ս7w;M�%�X���9 1�baǮ*�KҸ����Kh�	�5,'Y������p�B�DR��:"���S�q��Ma5�4�� iܨ?��h�5E��N;˕Nx�DF��@��@b~'��V24�9�Y`P�ء4���95�6��K0h�ؗ,����cіScՍ[¹3\�&::*RmQ�`\��<J:���c+v������f����<��Rd���g�mGb�c�k���EM�]j��!���&��s,���
IPL)�b�:u�ǞM���a"�i"�]��=� ?�kD�ۉ'p��k�2��%�VU�+$�?�|5#PКy���cWL���X*�:Ԃ�eb^��ޢ��4Y��xU�1����Ӄ��x�A��˼x�O�D�8��z
���*�Y|Y+��ɏD>R��\P�� g�T�Z�@��c�
���nG�E�����X�X&�+D������zc)V��<����T���%E|s8��m����+��I�L�f2��1Vԛ=�Jy-�$v�〮V����	aB����en��tYҸ��$�ƶ=�c��Y�fNLIp��(c j�K*enX�d�u� ���֐_�B�χ�cwc.�(�X��+p���j��+�X/��+��%��ޘ�~i�TDnq��VDz�A��Y�"���4��fRh�����U�2ˠ�y%�S#"frViوR��P��*��}�Y"�ݱ��ſV�Tgȡz���0�lܟoLeS�2l�����^ʬ��10P~3��:V��*�vb���.!Jy2*�g�&��()�R�\�������N���s0�\\<w�R&D��YeX��Xbx�w�+n	�fV2;����Y���q��7��k"�ۂTWDJn�!c)��/�z����%G,�5�c~3��-D3�B�
<cp�l�bWs��#WY2Q��;W��_=(�F��b�X��4�K3s�xV�?��+˒6�#L�>U�TFfǯUK�Iz��i�^
;=H�k�A��R2�Q"�1*��>r�T��&�-*�|�U�W��Ō ��*ZX��ZP�J���F�G?y�3"�ӓs��0�iO��6�v�g��Λ�� t_3#�ɛ������X�Sʔuc�Y�a���+pH�;����c<X��j�ʐ¤N[c�|�LyҎ�j�	���P��!}1��LeGw�E!*e�#���7U�8���ꔑN ��,���'�FVU�)֓2�㣃5^&��R-B�)��*���0�U��]�|�8�F��ϊ��i���vb�p�QJ����,��Ǽ��lyp�δXF������j9���P&Σ��9P><� �*��&��P��iN	�n+�dE��wm�Y3D�Le��x�7��0V_ܺ��MO.G��U�n.|� c����Tw��R0���i�w�O�߲�,�I���I���[�+��dqt�,�Zx��vL���}1�x�ْiF�P�Fe&R�Ze��a? 6�
������9��X���H��vA8�ߋ[��fWPI�
�7*�1�-���ž�����V���˟���4`�Y�uPX��a�%�%�"�T��@!M�xāM�����1�l�'L��z�z7�K���f�������KRs,Z��錹#~-�@o�rt���$��`\ќ�UH�(�"�c"	�ț�ͫkd]�d�v��Zr��6�w^wn%�)��
�sƦ:�<|JR�[@FrLl��6��	L�]_�qcS�a_���Z��n#��%�ɿt�V��q�
c錒���8᫹�g9Se򈳃d�d�L�
�l� }�H`�n�D��e\��� �%2I�S��drU�y7O�Ϧ0��2"�V�=���c�I~�cxŶ�����;2qû��L �Ǜ���+lrK5	$���A�Tc��A��1�x�t[]��.<���)m��� =1�H��UfJl�ɮ8cVDl܆`Կ�9w
�Z�U�
�����Az?�N�iZs����ptnmD���@i���2��_=�p�[�+̦Ei9��sj��4B���B1I��Ɍ����m�Rь��h�6l�1�5v/�o�pQ[��~,b$kY�ء�ZTϲ�W���T4jR���Tp�.�Qv_Ld�)�o���c[�#�Fb��QrR!�Qº�U�΋��X��M+C��J:v��J1�Qq!{�1*
��;7(&�~   nlG׿��;����� g�����3t��w�6��5\L��Һ�P�M3�c�N���^�ȿ�xb��)�gฦ����VY9E�,Q���VP��c �-쐼(䃔V��Z9���J�މ���@�O�8�#��X5�t�;�սo؟r�Kg�t�WuL�}��.���O/N��8fɎ��=Z�
���ivR� Q�ko4�NޘζB��*?wwolnHY;� ���%Q��k9f�2��B?��YC~�?!<J�0����o{��o�]��v^����^���4�7U���v�A�^����Į�ҚT��>�y|��ի)���0s��~����R�ٚ��as'!x#�Ibn|!Y{[��~}�����W ��Fu��z������!��I �w[�~���u�,]7�����2�~�t�M�Q��S�]U�˛��o�Ke��.���H���{����meI�_aT��O�`O-ǾsҤU4�k�ʂ���$�8���;�s��?~sZ�� �c�m�Λ�c�d�T�R>~H��m�����H@��<��?��� !��h�Q�O��������G����x��r#)��Z�;MD�"{�'�0��*Ƶ�O�vCH���� 8�Ǿ~���ʹ�Џ#BUO۞=�IǏ\,�h�⾟mrz>heq<�hĦ�К��x�}��������qj�O��G�� /����eEVHA�y�g矫�?˜�Mgj��i�f�s<8Q�E䬭v%���;��`�=~U�:?�H�Xv�?�9���� L��hxe�I$ ��O��� �=�wO_��Y��I�Ӗ�U�ہ+���K�8�'b?�{����Cy��Ʋ�������z��������V��3~�v��ݧ�� nG���6}Q�n����޽�O�-�gmcU�2��L�I��5��¶��Q+���Pw���i��?�:Ɲ* ����S���I+�s��Ə��J��6g�B	�%x����>ô�����=�j;Aԝ����Lu�m:ϯ�Γ�:�M�ֻ��hy���g9�#}w$S�z�7.�����Ƚ�RD���6���/Ÿ�h�hc@emF��+���d��E夑�H���1Uo-[q�M_�z������7��1�'w�W�PW��<*'�I��#�>�=����I���+���<��B{��'Zt�w��x��8�1��=�z���t�RyX�n�f�����Z&�r�G���V
ZGQ�C�Ά-�i���u!! 	-�EzM�K�U� ��`�{�"�Kc�&�}�[B]KK��X�-�q_���%Bg��jV�+/�V䃺=��'uO�����w���t~��h�y�.�ϻ9}��Pk�����tޑ�Ӫ�E�*r3����\K�?^Ͷ~��K�~�oE���u?p��z,Z�;�Av�'�(�+�~�
�f�(j�kī9iI ����Z��cխ��l�T�y&�����vz�,�;6�Uc{4l�+�X�Ӳy����G����gH�{I�f{�ޮ�u��޽��Hu�:+T���w+A�q��+�@u�l��h-�Y���Q6��ae�1���#�)��ku�wk]I��#��:�6�b�][`k��k�i� �Ta�m&��^�aFl�z����Y4:{KF
��3�+�h����3iu,v?l�w	��#�!s(`����q��N��������G����/��qӽͧW���?K�6?���i���T�2;�M�c�A�8U.r�Ҏ��5m�����KR�w����ӋK�'������ַ$��^2����V"Jd7Ԯ�u�Y�h�d��=����Kw��z�R���)If=�	Pw�p����n^�:k��w����{3�+؞�����];ҝ�=����_K:�n'JKR�&�l�	��8,xM7q�#N�� G����}��zźv.�QnkI�%�-�S�e�ϖf21i�8�hb�#�S���3��}vOQ��h��lI2��c�5Z�M%Ci������gg�a�C��/O�����;=�b����N�uGy���O܆^>�������|�-O9�诪f�V8�zx��1�e�����%~�uWp��ڕ���f�NA4�5����y<P*ƈOh?/Z2diY�i�Yz���`���.��z�ծ�Z���0A>`�0���<�J��a�EG
�d�q�O~���ꮢ����~������塛��9]1�t��}_K�`O���7T�j�#7�F<r�E�� `'�U�H�N��&��ZY��b�ڭ{6d}l+a� �ń2�G=����?�ѿ�m�I�B�Fݾ}2hk�Gl��fy �^�`R�����=�����ߌ�K���v��k���� L�r�=���J���[e��V��ҳuM#����,��Z��!l`��)y�:�	�ѽG�:�n�tϨqI��Lu�G�*���� -�ఒ#���� ��dR�Z�� �k=!�o`ud:�}�4�O$C2|��bh�X��|Ɇ9a��x�����~��ҽ��c��Of�cu�[��tu��n����A�䮩�Ryp�5*~WP��'�b���vc��%�ml�� �qnMŨ� Y�>�U�Q�75�ԥ�K;�fp�f0+�cWvh� �fȻp�������jh�@�hY�P�fH���v�Yj҆�:D�ƶp�Y@I'��42�_����ֽ�����|���/��j}+���B��z��:S_������+Q��ԅ�m	��ؕ�h}c[_�H�}ݫ�[oU��v�F3={�jس���<Ii<b�[�c�����wW�l_�[r��ӷ&���e�h-؎���vn`�f[ɕ 2@ͿW"^����ѳu?��{��V��^�=�_�>��GU�o���]��&��=�u���~�����M�2�����!\k��r1<q$����3�/N�Eԙt���P�JX�ŵ���Q�3�l7��B��&8�����������kP�3lD�5��<��\�h"�Y�����%��%a$���C3|Ą�j�Ob��}��u�Oi�_�=��~��o�zJ�t\��|��ɾ��G��3q5.�\lR��M$!��Z�4I�#���{C��94��Q@�����rdTa�]�h��{�'��d�mnX5�R�j��i���^5��01�2R����EU!I_@��&��_�:~ݠ�쮷���Zk�՚_s�I��Y��oz�O�����:����OM��qst]�5��p�=d�t˒*<kr��"����Pѱ�R	�ʄ,8h\v�By9hH�B���U��ļ)�"?�=+'pa��20~��?P�z���F�C�nS�s];���=�� ^g���Y��'O��^t>��U� �+?LI�Q)�9��$֫aV�T�Qy4�of�+#��=����3FI^����ӗ��ؒ���*�%H�2�t]����@�wqWG����۾�FL�����	㌶�����w��~0��Ӱ�i}��(��%����ͧ�MC2��}F����d�O��
��z3A���������I��}{m�zG���}O��l2������:�\�n����鮅���&��鞕�����O@�t�9�FE��rfYK&������KWX�D�����I��E��ϮG{L����B<�n�O?@��Gܒ��?ᙫ���G�7Um~OF��V�z��<X�^DA3_�:��,N��[0Yc��ϟ)ɰ��ͣS�e���I�U��O�'?o"{˽����euK�eS�|nÑ�n>����H��ff� �{��~�����kZY����L]Z޹�4�a��#�ppn�C�-��o��\k�|J�>V^>��+��x0��'�d3�� �s�]�a[i��Gߔ�����S�LH�Y��=<�
�������d�ۺ�錓I��4�Q2��*PV�(�wW�~U�#5�SFp����
�#=�b2.�-9Taa�<rć�#9 Ą�Ffo��&�!�*�*�:�U��&g�?1����S�/-�y"�'�r��;��sVK�]��*��f]A����Y�9a�(C�D��',\�?�)U?��~B� .Ô˱A
wc!*F�'|F8����C/ƭ<��蟚�x��g�`3*xBw$���FT֎Ԥ�_2V	g>%����O qP�2 L$��1��y�9W$�5P*�g'%�1
�ݐ�Y*�Ld�$h�3೵��� �,*_ŧ@�_��VwC��X�I�7���Q�%���J��މ<c�A��B�g0wb�D\\l���9�K��1Mg�ydIid���t�E%��a����\!%�'<�Je ��7G	j��UM9"� P��(���cdƬT틌�7�ǖ;��"Yysv����⁶>5f}�o��\qzN�),��3V�������݄P9#fX�ۀ�����PҊ����S2"�V�'��E��"���3 Wc	v�ҩ\�Z�-�k-���Y�Vd��շ��(wtVc(�ZJ(��Z�]��R25��H��mې����v]���l�O�c �I���aDc0W���A�����ܜ��2�=1�\�� Ӛ�3c�4d��n3������T?b��2��ffm�3�+:�{����ƍ��ؔs���8�cBʳ�<���oS!_�Y�#�[�@�ʪ�5��Ռp���K�)	� ׶5aɓ�c��̭P� nc���l�j2�n����c����DR�����1�+�vo���:x�vs��2����g9�3V��u��EBsR��i��s�Q�<3�Y���m�U&XcQ�ά��h6uu>,aUyJ W�r�)@�xu��%E]�2g���[�d���I�ф� �-YI�)i��k ���/<UW�G��W%�v2�
����"�hLX�<C�dc:#+G�d;M~��*���i2+�Dc��D֖�a�b�@���;\�Pї`�,b�D2wZ�x�4ǶD�㖕��1E���uF��|XȪ&s�%lܣP�xO�D��JL僫5U�;+m0@��\0��_lw���ʗ9/�[����,� l���1<m�1�͊��A@牴�s
we��I���9#�ࠖ0	%��͎Հ*�W.�_*qv���{����n� S�!f1����~U�c��J�H�W3�$�1]��U�eW�X�2eI7�'�rx����(h�Ld��Y�&G��0��,�[m��9�s�
!U�j��I�;�؂��-"F������Rl��S��IJ;ȌW*�\�D����X�N�F�ǩ8�,�4�LR��x�̟��*�FP���xң������7Lb���Uf� 
��$���e#c���&B�����-�ǹWʡZb����I�b���@RK1�4c�U�US���P�'Ǖ:	#����37��|����N������VC�"�H��x��˭�Y�M��>�� 8���cr\\z�8���>[;<�DV�7]�I���L�c.�"��G5k��\�gYU�EUׂ��(���܀�i�J���@�D���<�8��N�R|@'����}"��>�A$�ִ�>��$��٤�q��lX�T�%c<Vk�%�T�Ub��_�S�1��҇�~H�@B���C��1��|��-8���r���G���
"��#~ca�r>O���MdgKl����+YQ����x���۫nX��G(|�3��8��ro�)�jΠ��K�]h�J�ێ,a6��I�ɍ��R<NK-���&d �y3 ?�0V��&X�S%����b.�szRm.����]�o#���=1�Ƌe3R�Fy4o���䛳c�\�o:�M����*���"H�-:[���pwhE;�Ӳ+��ݶ~+��1q�c�(/KN�2
�h���A�F��tU��+��IoLe�p�h�<�O�P���<�6i�ݸ�!�l�@c�NN�@D�FU�*ӛ��b�
됶��%s����c��#�#Ӭf�;Q��z��b��	Y�*C�#��2�PY|���Rѭq��\�w��3�rC��c�o�ֱ��s��#��h������a��3LeVT���3U�h��i���˫ ux��o�����f1�N����T�x+�)埓��3�vo��2���q�	L�vɡ��h�� �x�Ԁ�Ob�K�F��g+H6�C:���0L��0��-�b�P~8���ǂ²���(*�Z�@T+-�R|v�A$����錇*�r�Xb���TȦNMr�,|eoɧ�#�0xQ�PIo��S�bgY5��#!�<VglWǮO"��%�F��<U�m&���c/�D&4!�+/��Z�W*	�������n��9/4���?��.�L����� ���į%��ADt�� ���i"&EU��E
�$�~�/%k~�<U������7
~�������I||UfI�Q��3I��{Я�0�q,�*��Rl8�Aͧ4�
xm2�	���,oR+�/5�g��R���J ���	N��!���'��7oLd��2o6���)�6Q{-$�ޒciE���A,v&[�`�����tb���X���Fg&�h�M\͌�%3K,�F2fʪ�`�F'��	�sĢ�Ѿ�.�����HI�����uv�g̚���o�q˱��Q�jd��3����@-6�e̐���3)����7�w�ʲ�K1�����+���i���B2O<������ ~*��_�ŤX�J`m�Q���9BJ�(+9�9{���H�;s*1�� V�Ȥ�'x�J��ʛ$���z�� '�Y;1$�Xï'4����X@�V5�m<����ZRJ8uP��n 1�rdϐ�u�i<zPG��W��v�ش�R��rnAJ��w��F{b�f2 ,�q������k
uec�*C3&S����[%yE�sL�|�JT�7�������~=�+�ȼAh��6�:��(�;�DM
y�,_����\ംj#�%��҃�f��U�ěw]�ي�0��qWW�]�m�U�)���~)o�2U�-��S����8�ι���J�^wת��9~>��,�i��3To�]1��S���π|����EQT��/bU�>7�� O����Y�%Ts���� �k�O�U��F��tEt� ���ˣzGSѳ5��Zucuf���s���t�n�N�F��|��UB����}�XF�ww2�,BT���.��Gk�ZR�Y��Ѹ*r�cT�I�v�$i)F^{��d��A w^Ld�e!��7�ok~���v뫻��۫0�ݳ��M]�\\a굍�����zm2��WMwF�͒~5���/�iZ�� �O��O��Ego*��H�� {RD�X��T�;Ov^)j�97bs1^�xQ��W� �e	���%H�9�=Y��gZ车��ܯ}o�oP��_�i��N��dbx;-�:�g���]���'Q��l9�G˦�t� ������ºz�h���G�$'��Xs��������?F�9�rh�H8�@~��>��H.x��@�I9�=���ζ׳z����]Ɜ�<�����:�6����f�[ff��T!�,�19" UH��VrUBrH�>�?���� �]%�H׃���q�ۏ�� �cӺ[P�Ңm�Q[Y��x��H�*l~Wr��b�:J� ����?`	<��/��?��J�^n+G���ǿ�_|�&��i�Q�h6>.�Wty1+��m�RN� ���r�ȥ�g,���<G����<�i�dv�����������)��F�ɛ�����\�e�%����%��ԑ���G�4t/B�	�$ 2�*�@�����y���j�����y�O �?����� ȺGo)�:����Yb����Dv��Z2��_��@'�����N�m":����a�q�?S��p=�?�[g�]I�)��Lkϡ�<� /ӟ����� G�OO�����qrd]��Z�Wa��b�S�3ğ^�&��T�[JԢ�bD<(`���?�B�x��<"�Ι<S]�$QFGq�<ه'�O����1:��ֺ���i�XcO;X�030��#&�3 �Ip�L�06�!ӵ��$�Z���1D��$�P���=qϿ�9��n��I��#�>�̅x^	��G���2�a�~��Wn����#��i�Z�Ca���=/�1z�����Z��#@��0����>>=56��>|癓��A!/m
[c��J�f��N��e�4���kN�Ğ*���"V1/���Y�R��`��Yjl���;*,6c?ٖ�Ey@!�*��v����wT�'�s��%�>��Ɨ�=%�ۺZ�7�<���q����=[]X��h���y���αʶ������g4e�Ui�Is�cE�gN7/NzO�� �B�ֿ�V���)Y�&��D5�7�S,�^���ױ���*_�[�B�]E��j�-q�@Vm2G����&��;�RNsQ[�'�?�/V���=s�s=C�m���w[�ޣ���cu��a�ڎ�֝��C�z{�8ѵ%�y�E�m�1<L�4�C��W�H:����Д
rj-�W����1�č��x�� i�Q2�� ��n���lA�ӃT7�/����c�s����@U�s�9N�;����p�>��^���z��{~�gi����i9��{��^�j�웷�9��г�����?���OA�2�}BX�/�4�qsS�m���m�Ӎ��:)��\�J�)�R�^�����#�O=��%}����RM�-P��² �}m������������uWh��$��8c�V��1Vg��2�#�ְS3�5=��2�GQ{��p�;߯h���۴����h����:SI�d�:f?O�&*C����⮙����"2��T��=���W��N�lkV�Q�t�N��Cf��b��<�Z�&MC�'v�U����l*���b�GM�@��>��qo

�N���Z����OMTyk� ��� ��D����p�JOm}��� p��^��ïv�R����vk�zw�]���e�C��gu�p1����j��1���Fg51&�i�5x?eF� V��r)�]ѡC^	I[p��'aC1�H#�$��Ĭ�������:փf�m�~)���0�~��e,�c ��M�Q����%�?h�����?۟fx��+u�n{o���Pw���M7OM.���,�0�ln�]%�wK�Ǒ,��ŦBD�v��k�?�];H��׌nY�Zrڽqi�-�����)唋2:�*$��cy;9�p��{� �oQ�:��G����؎�Z���TR�I<բ���
<|��2s+Gw:v�����u���7l}�{&�"v������3q���o��ιɧgNٗásE��7KY�������N��,ܔ�g�6�͝6xg[��#@a� u�3��ɒ#�~H�,��h������p�.�?��M�k�ԫM	�r{	5+(KΟ���"�L��'c�VE�1?I{����巸>�{e����q�ji=)���I�}1����4�����MSO�,��(�x$��ǜF��/��׎��u9�iKy�&��#���ՠ���@2�ӕ�7��26���k�؟E�eʋ�Y��:�0%� {$-4�>��$X���$�W�F{�a����?�_�� �N��^���L� ־���k4!�wG�^8�m����d�E���Llh�'���b�aƥ}^��Ǯ����n�h�#�6L0R�k�f��D��Q`AY�+��3�C,ݲJ"U�s�ۯ��/R7��e���;Z�
�Z�I<ej�gI��*�d�1pc�����r��j���hu?r��:�H�e���%׵���'{:W'��u�����\Ɔ((2���YK�A����X��R� ��^�|{hQ��*�Z��b敨i�+C$q�_5ײX�)��wt+,SC,`�?��u��5��.��d�R���j�u��ye�f��C�w�����+�������e�Mw�~޿O=7�}an��0:_�3{��=��,hf��N����(ϧ��z��1C�:>;���o�^�t;X���=���r+bD��+I� ��X��JÅ�j���L)�a�~ :�����綗j�U�岂��ڿ�GN��a�RZo�(J�&pC����V�^H뎱��N/Sk�q���i��V��n���s����~����.���1dOU�ud��1t��؅lj:��/5D�����*���*���Q�#�`y<��E*��P��_�̈́�0�i�?沈4��䓒�{����~�P�WCu��.��zߴ;�e�P���N��t�\8���=�ӵ=#�u��*Ox8�r��ͱ��k�~�f�L���m������`�+M�?T$�O�9ˮ�cU�aPI�ջG$�Я�� 	� ��(��o�p�����7��o�]?�}�� X���9Y����뚖���Mw*ö��<mK.��.��=�gK���Y��iW3O�#�1
5x~]�g�y�繛������ y'��,@��/l�y�W�@�
?_��I>Ϯ� I'��\�2z��z,���T�>�vy ������]��?�F�4�S� ����SU͕2n,��f���K7$�#%��A<� C�Go�#���K0�����'�{A���$���;?���;Uَ�tgo�����S�X��G�������k#N�s��G�s��֔˝��W:YU/[�˔%,W��ٌ!����99nc�����7�����%}�,�keܙ�s� T!�Uq�8en>���I=�v�{��_���kB��+��:��\\.�������jX�s�*j}1����ɓ�긞Pr�h�z�Z�wSגt��h}}|��pĨ"sё��;I��E֭}1�n"� ��v4NC#D�z�4��zwd4|^��ƥ�՝u������B����W�5��3Һ���5!�'��In�ȝ��M1芞�]�p/��E1 )\rݧ�C�TϜ���z�v/�TrH^
���럷�8�7�?Ժ���w� 
��ٸ��:'���|��TմΤ���|�;Һ�]p����A>!٘oo���% �p>��U�ߓ��U�&F$��� >O�8κη�:U�õ2q1ڏ�����c�`�h̠�-�h����,���G�c��cȥ->ynӡD����r
>XʲS%TV�l���w�Ĉ�0ѷ�V�jb�M����k�cz������2#�I���h�Lh�1^��p��,��F�l���1��>E-k�j�((��$�@�����J����&D`Oь�mXfR��YN<`�Ã4T��gy�ӓ1bGٙT2g��{��/��9�,�H��c̛�J��}׊��(����Cȑ's3��z��9g��ʣ��mj��ށ���'UX�6J��;d+�c��㫿./:95BADZIF5�ɸ	�Cq��|��ly�*>4g3I�T:��1\��)4Y��,doh���C�64���Sz��C���x��U��ȱ����ec.D
�����F�m�b�h�E�7޳)�0ك�c���;��X��u�?�E\���!�n-@�4�nfHVa"<i�A��bR^o�Ʋ��W�F��pt��8*D
Wn$�c �JU���*e%�Hɐ��{�$<>�v^ ��eW�24�9�%����)�f|t��J�<@P&�ۊ��b�f2���j³����3�W1�^��T��`�Q�W<�7"���TǌYC孝Q���txU���B��/��@6�w�'�|@1fj�ue񌻻�"(��к kYf�$X�q,W�]Ճ(`�����9f��T�uɉ���"3ƚ/N�
6��T�'(ڍ��Id�_x#7�E�$�-0���ͷa�9*��Y�u���\��/�L�b*~9���1cP���y����,�d3�D��bk'.�4^Sv���c�ș決
Yi�Z�*�k���t)_6���<{�q��ec#�UhS�-P��\oE��-�4���I���1�w��y^SEjK�..N?&I�H���g�UR��P�U�(���&�/v��뒫\7Z��?fr)V}��F�p
�[�:Q�v�5y�C�US�d�Ĩ�(X;M�)���ݛ���G�m�rq+�껛�h���w��n�X�P|bn��^f���q	��~0*|%T� >U�M�1�Lud�mĂcS�,�j�	�13�N,fHD<�<d1�/��j�%VV�$���V�f�[~A<P�v�y����7��'a8�tw�Nn�D.�����\�5��!�8&g��1^�4;�LLw�z�w��$iF�2�
$���b�^$�c	&*�8�T�ԕk��J/3��G|}����hhFͺ���+�ˊ��0�Ia6�ȜS�m����;�&fA��5a&�k0d� ���2�7��	�ƿ�oo�n�c`�X%))<jY�Z��2;!y|�_�[��ɻ5����F��]KyS'|bl��s�Uv.	��H�&�-u��1)"&�_ �ȼ|��)��@c"��yr�תI�}������qiS&�B�`Y��t�������;#%����fT%���� �����쾘��QSC�I�&aR�1�NesPM��Z��ʣ�`8��I���&D�5h_bl�+��XKlZ#`�J��� oT*�^P��V'��<�L��0t���2�df�8�.�iĭ<i���z��Ī2��Y�?2A�}��)e������Ȟ<ď�������IX�U]�@�"���"���=�]�������@��)M��<	ߏ6p�0���k_�d%�&��LH���1�Gv��`�Y����Z�e���/�h����-E�~	�	�~�����<�*�����K�VN$�P�EM����@���f1i�6�B�3򖟒g�Er9�ќc�
�� ��"�w'�!X�(bbO�0Rx��
&/��q5z�~�C�
;��/�WD<UZ$���l�ɋ�R�V��1o<f�H�Ď!~W�_�?�������2
� ��f���;3��r&��,di�*�'j2Ml��rvQ:��)����� ҟ<
��c�ƜY���Lv��jЛXV�� ����\�R�d�F/Tf�=9�V���
�Ⓜ�� rZ��3f2�<kR�3� �]��ߓ7"X1	��5y�E%������2s8�W�a��ew����%ri�3W�2Wz����T��by!�qŠ�����_UI��"�J��YN����<�"�i/�uVk���<u?{#nJ��T*eP�ޘ�]8�������ǎ� �u��o�����$d�E�
d2ٲk$|U�Dk8:$����Pf��>�eb�nm��<�/|H��z-<e�4��c5 7��;Ld�W��X(�4b�v"SY��Vg�QdYM��C��g��>c���l)$f	� q ��I۟����c'��T��C	I�f��aZ+yc̩w�5!'�B�,e�d�u��!%{d����J�c��D$���Ŷ]���9�½RT)��?�ڱ����b�x&����� �8c
����VV�kO%&���s$(^n�t�����z��5Z�Uw�%- k|g�8�˹�V�8s9L.�ޘĥ	�C5$�c2�ς���b�D�� �ۻҟ!Q@)�zb�W��&rf�������'�~ ��N�zc 5�ߕ�3��m&�������z2���!��y��� �&���$��e�f��A	�w�*�b����Yx/�Hp�錐�I�;b�1wvc%*��,wf7q��Y��wkyG؂�Bh�jPd/0.��?l�uaZy'��,~=1�l�_9`������S1�X�E����X�UT>��-��ĶV3�a�zx2̍�M�ԥ)J�x�
Xŭ����Ǹ�����a*O*�'�D��) q*�Ēx��1q���W�Ix�9`ϕ�_-��
)�U����X�H�S(cq	���y��/�K<W�����Μ������x�c��O$d.��Tc��NU*g�]M"l����(Y���d�c�h_+&G�%�J���T�Z�B�[$��w�?�' �M�]��k$~K+��K��o|�j�mQ.C��.Qx�����b�̓J�e� q��K����b���E�V��!�vV0�C&��D��4UW�q�����/��r^'�/
د�c�'�Jh�J#sP�6���I���,柴����?�k����l�c�fhJ�.&,#���F�.4\ZUg� q}��$ I�3���^���2���h������Z��#>���]{[��lCP[�q��2���$G�2\�!�d:v�-��ZR<z���[��#v�UJc�{߅=�I�9�$?4!�F�I/r�!y?�@�� ¤�g��U�eٟp}U�uҙ98�W��ƕ��ȍ:C;/Oֳtl\�c	Z���A�:�ѭt��_G�jmm��֫cMi"��G	�2�*�%>�䟪�ø���<���OVYⲫ,e�Oh,�r Yc �(����=PIs��s~ǻ���[վ���?���Mo��њ^{ә��f�L�]D�F��u^n53�-2��&;�꺖�fo���1S���|	�!�n�b�Ox��߾/�iU�b��H;d� �� 8d�^@���v��#0w=�utR�#-/L�oi�֖gN����s�|��c���z�C���u5|e��jl�y2bc��V~�.=�G��Yi߸� *�'�x���O9�Z8)~����� �p��r?�?�����a|�c�J���F���6d ��I����?�7��T�J���}~G��?ZX�(�������˞�К�����*5�2K#�;H?���(��� ������,G%V2��~��?˃�r�>�r~ވ���O�d��K'E�u!��dOt|�ݱ�EIqG�l�3���s�}|�16���~uc�ҐrG����ߠsλd�fO�g�rA�~	�9�� 3�ɝ?Ӵ�u\��gQ1�J�"�*�U4�\��%�c�7��_)�� H��Y ������q��q�T���w<���߿��� �h��q�ۯos�Ĉ}�aTW,ȸ�<�P�ȹ�̛����ۃAI~ZmYa�}8n=�<~�P~��$��JFd��n��|\���^�F��>�����N���^5��]���G�v{U��b~7�5�.ͩkjU ]^�r���CwrA@�w�������]�����m>�]���r9u�y��3���L�jz�m�]��Su?K�:U��Z�&������>n��|���rOĆ=ml�(%&��4��������2iF�� m�rĐU�����*��� 1$���ˡhqE�D޳�H�a����4Ĉ�bù�h`�ʿ�FoG�_c��힋�����������֙�&������{o�i�u8�_ٮ�3m5�FF��z������Ҕ*�p�	5i�S�����j�*���[M՝8�>١� mPc�V)���&>�����ܔݫ�Wd�H��ػZ6����1K�R���P�g����wP�#�;��W�.�wǸ�Mڞ�e��C���������t����~���t^^^n�����r�.��g�:S:���N�W��^���|�Qv���jORDRV���4[���~CS�5��~���DճY�HN�Vf,���=���h���wk=�5
�R�=��S�G��E�K�L�X|M,qGh��{�k��O���tM{���X�m{�:GLw���]� ���8~�{1ԙt�4^����L7Z�ji����㮩�h��ӧ]=�]#�	��ۨi��L㔸�jkZ}m��D�u�yI�ä���˓x�%}uJ���_F�v�r�x��Rv-��jH待����V�yٛ��}��Gw����+ٷl}��Y������'I�1N�j�e�Υ��������wQ�+�u�U>��)mX��p��q�tf�)i�[C⏢�.赼w��7��*��v�H��*}�td�eE� ^�^e]��A�k�R�mE��v�퍱]X�!�$I|��^�� ��+�HDa*T�*Ι��{"��ϿQދ�	����T\��z�ۯ��t��^���w}s���2�|�M��z�ZQ�� �����l_���t�_R)O�u	�==Ml�+��z�G�F� 1/^x��pbc$kJ��S�?�t�+�&ΐ��~*�MY��񇒲���#���WI�p�J�`�#�t����~�_�?n{����s��;���p~�:�F��OF���MO#F�S��y�L���8�l��9���l��:s���|!ӏ��X��w6ߖ-;O�bu��ߊH[�,x��a2�
�*�<����?�Į�� f�E��5�ś��סFX�7lq��K��N����L����?����Ϸm:O�1е>�[�#иy=��p�Q��+R�����'U����Jk��$�<�KU�k��~���ӵ}akP����w��� �"7qS=%�4���v#px��MF���t����pX�#+������3K]n�(�]{���]���߮����� g_������t}��?�}�=��/x5>�k��nu]3O�3]�������FfvP_�ϋ,�ȥm��૧� 6+u��[��փwf���C�l�2=�ׁ O�3�(�9�3�YP[vgņ��f[�&�:4�:
VH,��R�aYE)�ʁ��n�yU�vE�H�F������B:P{���^��Q쟶q�{���Zֿ�wK��A='#?�uF���#V�-�vH���V���q�9�.��O��:���2n���WN��R�M�ܳ+4���H�L@�	H`'r㺿Ww����?ӫ��[H�_���jjլB��׉D1ƭnhBD9fp$�~�dx}����9{��-����Q�N����ܝ���Z�-/'�5-fo�-2��v7M��.��t�
�da���&�����?�9���j�5��*x,�<uZ��Y�D��GnI]D���w�y_���	sqG����m\�o�-iR�	�2xZ����Tf*$��W w��O�����_��Ogݝ����r��}ܛ�MНe���:f�]�j�7
�P��Z��8�j"�<�L�}�/�7�ni�7uyzuG_G�h�|�l��WH��Yx�&�x�,�1�2�� ��/Fw6�����{�A�(%��J��MRͷ�)� Z�F�<���G,�8p���~�o������� �N��Dtu��O�;]��Vu�_�fl���mZ-N�uv&;�r�Z8��vw������:�OM�֡gJ�%�J�i]a�l�rU"2EJ�8*�$�H I�`
���'Z�tij=B�WW֌�[uP�)An>�)��j�ߺy"�U�x"_��\�~�=_ۻt��=yӝt5�ެ�z籺��-��X�&��t�_+S^�˦&���GLu����))kI�J�P�wi�
�xX$��$ts�w�T+�<rdy�ؾ|� �z��O~A�ʎ��:rC���/$s����}��<:Ƿ]�^��_��=߭k[�입�ZgLw[3�l֝c�5[��o�d^Y��&6�lz���)p��/�*j]�}ֳ�ۄ�H<�ah���j��|�H%Kv��R�e�@J�����x��p��d)��s�}O���~���ݗ��o|]/��)���v�O}����38��Q���v��?��:�_���5��^�y���,�(�ʠw�D� �J����8B��x^RK�'�x����^�=�{r��Խ+���+�o��ԸxZ���WS�Wl���G�twԤ:�^L٧-Jح|a��F�P�:v�,�盘"Ew�'�p�v� ��O����,aQ�3���B�X�9c� Q���+n�t?|u.�����Դ.��v�OM
iq�i鍕xch9Ԛ�u�
�U��ͥ�qF;��Z�>����h,-kj���݅��xW�.{���i!f_�A x$���or��t�y��VNo$q�(��ʳg*:ϴ]K����W�������dj}��'G�����3�,�|]CF���we�dt���|�����K��r)+eMgX푭�%2s�H1�Ҳ��!��'��nr�t?v���y�0>�+pX9�<��f;�us��G����Ei�O���	����С�O$�W׵�|޳�A���5=N���X���V��g2#H�Iq��<z }+�珿��.��@��4���������k�T鉗s��� 	+�ܖ��;>��3��@�׽y���G�3�X��~9���,�~0M�sL{d����u�(i!��P�����Qn&X#r8������� �<cp�=�����c;a��|�R؛��;�E8(��E��<�U��[��k*O#��2�%{��F@�\��>u��?��? �r�2r�7k�5�J��I���x�J��!� +�s�59Ld��si:XR�tȴû��*c,��6[[�* �Co���ŉ#֔��y9�5D�1��Kr�*�h���2�錨8�dΒCkņN>,���P�%�E;.ܝA +2у�1����I)���&�fUe>g�:��B�����1S����2�q)�e�e�Oˎ��r8���S�/����7rX6�2	��q+�U�"���vu�K���\��._��c��a��+���˦R��PZ��ˠ���y���P_}��,d\������#��db���J:�eWE��)I�W�ٌ�i��E%,�SF����M��@� (P���ucq�YR�|O<*���\%<lܖѪ��Y���+�e�C"tBο��*��t(����ˎ@���P��43�L����60V���&�Ƶgj	�h��� �����}1�lZ:=�l�ux�+v��]��%��M�O����c	�W��ihY�%�<e㪊c��䥙���x�@�c,Uezd҉�3�����[��n���y����g�}L`��:�W����z%"C�$�äd�f�<�U���1�*2�EᎋƔ�2�2���m�	W����w�n	��4�K�&����]!i[2UX���
Ա���?m�G՘��~l���7��*����92�v��_��hG��lZ�R��h��e������Y�����V,����X����+�Kic� ��p�I�v�Lvj~+&D�ʴ.��eWw�GL�;2ѳ-�{%&ғc�A/����N��N�)p7f0O1�LV��Fʶ���-rd��MnAP�O$,8��,b'��Y�CɓJQ����o���fk�%QMK8��5Q�'�-GJ��d����TJ!,�M�IF���~�X�y�.>�#�N"N��	�*�sG�_��eFc
Ù����9fPfJ����
�P���%��Тzci�����{.=x*IgJ$ �O+ό����@��H��v4ac@'���$ �B�^s�-T��g3c�rB1�:Q������|�L��.l�M�*����a��� (@׿�������G-lKx�,�|��X*)�W}�)(�Rr�]�p��W̱˴Z�nJ۷�x�AM��H,wVU��c	L\B��B�O$Xͧ�G_�ي�T���|��X��`�ǥ�u���
N��$�:�ԞT@���;=@�H�j������m0�����3X#�ɘ!N��`�{>�_�	����/�4� �y�/M�h����tc'dz��jS���|��'䗌�X��,K(�3��M��P��c0���cv�X�C�8���+����Ld����*M��Y��Ex��Ex���/�uU?����Ӆf��i&E��$%�:�{�������|�]��V2N,�X�!�l��x�Ճ;eI��x��CnK��,��g;J�/8uR�S+9�J�L�E�y&�p1�B��0�:S'�Ch�#��9�L�͂����ʠ�`�B������O�t��3C"FSp��+��:�����Ō�|����?�V��I��Kg����o��O'Q錨��H���V�8�ǒy%�d�V�N��Af�p9��cNl�fIp��ƹ5sU�m;ދ7 7�OuI��� f1UvƑ��ä�閗��$�4G��?=�|�UF�l���D��"-�T@�(������%Vv(��9p���B@ђj�4�9c8QT�LQ�-����{ C6�a�m&�g7I ��I(|v��F�6�8qeQ�f1�3#��ơ���*�6o/ԝ��I�>��zcA�uE(c��)e�[URV���D
;?�
�t%CFH�&L�/<��A�Lx̶a�(��T����*X��cL�r����ź��*W�l��f/�x�Ͻ%2�;���+��]��d�96@+U�1�Q�	�GrǦ0jw�\^u�?���)�!�>��F}���b	�x�c��lg��i4�r���;aҋEǠ���Z�v%O�p����A�(l�4#)���YT<j�7�iQ�*�U�͑G]������)�?D��h����j�Q	0HP�'����3�$���r�SEi��"�<8�mL���NS4nAB��rG�07K�Q�.3�4�-��ˍI��JJ��O�U$��Bl�G&c��Jf�)i�]B����*���R�W<�N��H��?�X���#6qD>aA��v�|K*�@���7?�43���cyF�g���*�P�yK�-�t]��G�� �k�C0� �ٯ8��$���.�h�L�j��*�Ń�#��D2VF Q��yTl|�����<-GY6="嗓�G���zc p貔����UyR�����e6`i�F.�:8 ϶��
��M��(�#���Lɑddm�|͸�������O�~ݛy��_�0�M�ӡ���-�=�T4�$�,dU�G�1���4��1n3^)�V*M%���YB��wQE`�?��g7{^�u�4L�<�����|��x��k�e���=1���**$q��]j")I�
��BJĲ�m̓q-CňA�+ѸJAgT�d�I\Y(r���e��"MҜP*�ŏLe_���3%���RbKV&ߓ�i�H.�����a�1����4�<���y�)�U�$��d�}���|�Ld$���"�e	���m��lw���2�@t>F<�UK�!��ز���r9���Լ+A��De�9�����y1�&�sE�d&��c+T���Z!Ȫ`2���o���\\y�:c"����(�]����N\�E�&��Lc�e8�%��5�^�Ol�{�!%j��	c�*��
�1�`&&�b��⒬,���ũ�j�� ����P�2�H�Ys��k�c��)�UJ��y&jHB	_.˰c�Y�c�r��*���I��Ũ���k�#) �őO�1a�7ɫ�˳�+�^�n��^)��lZ<�Pس;�vTEd����;w}_�y�z>F���M��&3du�VH��w�ӌ���:�Z�Y�8X�� #"�K�v��Y�,�j���xD���>�~O��jP5���� 嘁�j���_�x��w��RG�2:+��.{Uн�=��"����WR���Qfu����?�gm�;b���R�idT�]:z�#����'p��ѡf��tfg�	G�/k�$5���b	!T2~�c����'p�Gּ�I�00��o��}�v7������to����\|���̽/Iҧ�.yT�z�J�ѻ{��m7���������8j�A^��i\J�\��8!�倩n�'ނ���Ε�?V�f��b%1�Ty�K�������>�s�]��Gm��tnN�xl~�w�m��[��}_�z_3/Ml,U�is�東oZ^}C��\��5��qcFS�u�m�4�3�[�׻��]��b����*~���\g�i)�읦wu!A�T��}L������sL��U����k�u���>���Z�}�SS��?�dgg�]��)���Y�u@ [��j@Q�?C�<�������\���������� � >�=+�Ƽ_#�0����%Fb���$�6�r���v����M5VIye$����������b8��-ґ��<~��'� |��D�ĭ5h�m,]�ʙ�Pn��2���7�q������iHG���y�
O����?�2U���� �[����㞗1�=VZM3ǔl;� ָ��ڄ���a)�VD���� tvu�n�4wT��Ǥ���IPx�������X���~ϣ��kH�~}�y�Gۑ��� x��{���\�6�������0�&�H�+Λ-j�`�x;
Q�����z��Z�~���kS��^A � [�\��-򴺜����ւ1�aϿ�����>��2F����\ޜ��1��2)��[i��T%0u�s�ŀ#�yN.��qY��j�5];V�{���ᇦF ��H>���񒆣BO��@��N��;~���=���n}�3�uT���r��	�&��^�u8^C2��qC+�b�Jq����ku��46�9�e�$�?P?�8��� |�MGN��Z������0`���~y�f�t������;S����~�uszs[��;\����.�����'].n���l�\���Xb�S5�Nf,���j�ޓ[�n�ڛNmR(u
�H��s֐;,A�_��y"��:����:��nǤ��K��M~r)���ʰO/,�?|~���2�>���oo^�:�R���]/�/b]���,=#/��=ԙ]Q�ú�qΒ����f������6Y�+���[T����MG(���O����=���nSù�Šj�E-UL�x~ƴٵ���3is�Zz����<�l�{��Z��ݝB�#�[n΃����N䖧� X��������1�3��"k���Y�����޸���u7T�PK��m;�=Eк�Ma�`j�_��}S���1;I���_�S��I�b|0:���+�F��V�ڥSL"����-G��/,��'��\n
�j��,��Mz�\v�V�[O���� ��Z��i�MF	�-G斪WQ�I3��r��/wS4���l��/�ga{������g�K݇w��+N���,㇬����G�r}��W&�Z�_Z�)���:fv%rw��;s�[O����ɥE�{QҪ
��;�u��.�bܞ���,:}qcR����\�a���Y�e���tڶmWq^����Q�Ի���R�fmN�,��di�'� 3��4[Q�o�������t������z7M�B��-��\�����vJ`jX�J[��p�i�����ѼPt�ݡ�/�?�2_�3���ck�7Ѥ��جڅPlC%{U�)5��3Ak�-�i �M�Ds�:{�.��:�>�췠4��R�b&��-yP0�����E�ݒ1+�z\���+�.��/Lv{�����ֻ����;���}7���?U;�S��WV�S�̮�։�)2+I�}�3:�CWV��]*����V�� >"(��U�N��f,I��Y���ސ�ɵ_Q�$�`���*� /����ho�B�~ٻ}Y�/J�g������ �Α�{���kZgNv�}���>��}N���{:����Þ=�l̲A�>���n=�?R�������Ι�t/g�m˨��\�vW�f�;�pV�䕕��JG��r��� $��[�{������Ӧ��^�|�j���h����4k��O+4�XI"�)����7�����~��Os��u�B{��wqz3;��s�=B�uu-79��OR�T���<�@����ľt��N��������%���u]�3ǧj:m�$�=F��)a�r�3F��RA,S,�vW���� ��n��ݩ����r�Oj��c}6Yf�)��VX�X�e�1	�o��V��/���]i���/鬺?yt@�/M�uW�n��>���X~Y�Өtnݜl}I�ؑ�)�<���$�M��{{B�"�:�,�mw_
}�F�;Qcig`�C#��x q�m_�I�V��K�����.#,�-ƫ!q��$��r�?�@�7`H/�����~K�7�_�g�=�ջ��U뎋�'`4M7	t����t��~V~���ӹ�"�"�f2���j-����}��馍��M��2^�<�a��-hbI.<�$��哻�q(�ҿ��k�r��\޺�u�kYJե��J���-
��Gfi�b*"�b{�Y%fc�z;�;U����I�������t�ns������k#�tK#��h:�q��1��tl�c[g�ΆLi/YN:���VEO�}R����V�h�]��-S�2�Yk�Ҫ���|.�RH�BF?�O�}c�K=F�ν6����<���ڗhY�(�$��w J#s�d�5x��h�����7LiYڿ������}���O����yzK�:����'=铪׶��<}?V���Cn�Uf��V,�ÿÿC�)�����Ϲ�p>A&Xj�x��o�:�
�O��QL>��Sݒ�����Y��_[���8 ܟ�,���R��p���K%~�� ��nd�އRw�R�~���.�Ǹ}M���w��X��]sT�^��Q�T���I��f����P�*��5��P�=GSV�J��i���QQK�4`$���r�{{��;�̆u��vli�a65y�{��Mʡ�ܝ�N�^�1(X�Us�{z�Ϡ��ҵ��{��c��SEյk{���sI�Gj}3��F3uGs4~��7CfDǞ�����2������t��I,�F�v�嚬�~�'C�! ���DÏ�`fEVޡF��B�=�āa #�X�5�$����p׿^�}��t�[W�_Jk�Wj��x]��{�~��Y�b����� �0�Z&r)Ȕz�Y\��hЦ���/kbU|������?[��*�Xq���'�����e�a�%0,m��}' ��h'����U>Ǽ���O��{�{������l;'��յ^�u_�j���ޣ����n��ur�]C���v}k5_S�$�H��Ɲ��x��������$�9$�� Κ{
f�}������ �9�~�ײ��~���a{_���I����Zfn���R����un��4�w3�;����KL� L�/'8�g��\q��21Q"�����%���f#ߏ���^]H p̬r
�W-0�>y�M*;��p$����.P�{�i v��s�:����H�7�.��='���SQ��?�2���.��'k��X��f0r���L�Q��
��]����$$�	�*��y�K+�fB;�vv�$���\���i3�����UW�U}s���8c�@�8���ή�{1�GB鞤���p�'Q�&���5�2�gJk�zu\�Lu&���r4�6D�X���\����8n�U��?�S���t���Ӻ��C{H��߆>���/����fn��|��W;,��Z��{ej:�[�O�����L��;}ݘ�����]i;�d_\}���.���x���m�ʑ��2Ec�u�mٕ$)ο�� o���n6`6�q��t崡�߮@�?��󘟏����?�甖F���G3�C��Ȏ|��x�??�A��Wm1R��C�9�z� �����3�7[D�>�� _��>����۹w��f��M#�)lJ�66N$5�E�Y0q�"^K� ���ei�c�mo����]\�ԍ��4_2V���^hܥ�����ik�1�C�9 +"0��u�{���G���ٚ��<��(,C*y*ه�H"�	�Ieb�J�%�ta�vw�;��k���&�u6^�:6rO �|�O��4e��A�$�,]U�T�;	lj�{�z�;I^.�Ր1MK4�������ܼQ�� ���C�m't4{tLU,KΝi�� �k�B������*O+z̵�1W��Z]Z������q\PܘMU�-yH�V���G�x��?|۠y ��� ��������oh/���#���kUS�7�Na����c����.$�H��"M6�Uǔ�!�E�ր݈/V�W���*�.�
qϕ�$�:x�-��X�#���ud�*��tQȆٶ`�*�V�����9����� o@��7�*���c'���k��J�s$��j)��<n�I�H
^�U1�����eIA'?:��#%�or���cy�m�,6a�2D�KF	X�G�^��r6ʫ�
9YW���2�]3n�`�qD��Z�c�s4Id��y�p`S�������ډJ�yC"���Aᩜ��S�6A���R��c"��@J���PG%���y
K�K͔	
,>���#�k1[7���h-J1�3dT5 
��@S�c�`�Mӣ5�ds�>���g�NI�Yȿ�}h� �8�b���v2��^J0���I����3��P(w��(꼋��1����\G�:~=E�/���x��U�
�1P���e�d��Bt�L�+r��*̎+=��EM��O�錋�ɞ�(/���"Lc<[9 �@��~EYU�6���eV2O*E�t������\IkG�R����lW�eQŌ�CUm���B�V(����i�g�'�]\&�6����|�s��JP��!��J=�6Yx�1q��B^�����vٌ:�#��uuA5��`��S�38�͐�&�K�?oLa]O�eRB�<�5j�Sl�����.�E�� �n`w�*�?�<9*�O���%)[� ���6e�����/�1?_�]���oƔ��T�J|��T�� �J�Vf1_t8�i
��e�!I3�F.խ��A�@��1n;�0�6��Y
��%�(�{G!UC"=v���|���s�o�Y�RŹ���h�!M<y,�4��(�h�,�/�m��Tcpg+-d&�w�[��j
"�S��2��]P(�fͽ1��2�X��0IT��W�J���L�h�lY�ۈ3v�� o�2CcR6<h3+��8�^	��"^$�]ܨ'�
 �����	V*�\tJMw4[�b4gy;^�Z!�3^�s��vT
����� �}���5��T��<N�i��J�	��c%d��	4�?��.ɐT�˥W�7*��b�@��	$/�\����%�����I�� K,��v��25�%8��)|b1h��5e}��f�f�ق���x�0�|d�FD`!��68��x\������KU,X03�31��*���	��||�%U^|qER'��$��umՔ1���n��o3��0vu9v����G&*��؏��a���J��ȕ��ț4	�����i��ʧ �]R�e,� �\�a@��j�z�R�ZP�68B���Z�A>��..�����O��1��$�@�������w� �c�=|V>Y�%|w�kEg�8j.��"I����(Y�ح��D'�
b�]�*:3-]��&`T�p�<Gt��H(��Jd�}�pm˙c+��ݚ<�J��c(�j�
МQ|a����O*#���i�ṃ"]��Z��5O%E��
HU�ٲp��r6v���T�܆0+���0��/_����o4v�fm��M��.D"��X�m�^S�x&,��Y�L����.	����	�+��0mZ��Vl���iX�U2�Le��G�*����b�)dZd�eBI��E����DZ3�V�6�6���$�P���W�E�'�<2ɝ%����yn�Ncg��7Vc�c&H!��L��,eP�bY]Ձ ��R�fJT�=�,dY�~?�C�V�ܸtj��R�4�5�a[c�\�c<v�[ƙyU�a4�KRc1�N�9�ʤQ�b�zc���P�Z.�_���m,��<�aYm�+�UX+34��.$�2�(T�`��"]��^��(���3;￦08�껽$�h��2K:���a�J'?��9�@>���FNCdR�>Tj*dN D��T��i�u�)�\�� .Ic+.Uld�� ��J�Qf��ZPd"�|@���T��e�b�S�� ���/��m����9��4�:Py�/UUVeUm���)��_3�Ee�.;3���-��_�f���I����2Q��"Z|�%�9͛�m�ݘ�>I?>��lA��g��ڻ�+h�X�d5�j����Q�:l�M��a	�k��r�ZYq
�K�l6VEF��9�T�Dd�>8X�����q)+�/a�/::�G'�����_LcW]��l"Am:B��y�jx�i�զ'�SvZ���^3�3. ��#�UÐ�/F��y��#��7�*89*G�1��J0��J�լb%���4�@K7��)�[b�Y?�=1����(�ȥ�N�"�uV�(U8`�*��s�a�U��Ƕ;a���c��N�h���k1UP%�̰P��Hŕ��_Ґ��Kd޳iO��� ���M8�� �����P�b�ȤeP�9�eVjd<��fr�9D!�Q8��dc~�U1�3<E�� �qf3�K)��ƲI�dZ��� �XƁ�^I��R��2���9��L��n(O	�<6g�c�O�b)�?"7İ97^
c���TY�<\:��@ ����9���'i�#�.E8���P<ԧ>e�[�2�yrv0VȞ=(j>B@RYa��BF���f>D��s �c*r�s?Q��儗
���G��R��[��P�>��2���P�ɶ-2lII����|�wF*���C��C%�L��vz*�֯'��࢟�1]�*Q����=1�č.W?��93�1�2&�� ݘY����(�!�`�ь���9)�P�H�X�%8�őr*mu�\��+|ېٌ�'K����S#�j6+c��ڠ�1�Jt!K�l
`'�:ݠʠ6@��ƶ�lj�p������7܉!H!C]�C��9���ɣVkiN&k[7*7
�X!]�f �ܶ`
B�f��..'����

�KЀ҈*y�6 ��x��6fWn{��e�3�����d6?�t��lV��£�rge�3���-��t�H�� �ϸ�2��Q��{ {�=�s�I0u-E�?�}/W�Gc�វ劣�_�]D���7�z�H\z7�7���&N6��Mr�� +0YR��]K���9̮8h�EC돭RHX��3�ܰ�[�<���+�v�#+��<��;$���ݟܿo���Wu4�qV�k�wϷ]k�����j�:V'^��-�}>��}�"gL�n�Ǯ1�uӆ���l8�R+\����u��v�{�Zp�`�)@t��w���83�x�%�.3�ӵ���U*��{�YRD<2/=�zo��A��]ގ`��{���-+�qzg�:E�VgL���:S��nt}B�ɶ����EPuE[(�5\�H�ˋ���N�4�8��P8�?H� �bI��BAB�y�r���<p=�׸&2dD�(�~2��F(Ϲ*�v�  ������RxE�O^�� ���2��˾��v�ƞ;_O����yp��w<��HR�,� ��^�����"+�)���G�_��Ϲh̩�J��>���� �#tχ
��5l���n1_q,b�p�2@�o��?�o^�k�G�z�a�]y����ײG��yV�S2U��6�ڐ9RG�9�?���LSX�[�2��җ���<x�>[f\���I�%��$�7>�#�ux�d �\��y�I�\g�߭(/̇�W�$����s&ϦO�i4��uBcթ�Բ�͐[��Ś?�u�������E��͢�jD���# r��������px�z�x��I���=Ž1 ����y�� �[ٰ��d�Ư�P.FFfJ^�փR�s��0�>^�	�X�E��@��-[�N�SZ��<z�J��{��V�P?��ǣ��h�֋�CQ���3/�I =���H}r.=����{��=������n��z�^A�->Y:_�];��KO9o���3���L��'?���T�vF���v�=�^���-�w�Oz�`��ܼ��@�AbO���wr�v8䵨5魼U��^	f�ilȱF%^I.�=/�~�:m��wp=��^7�N�{E�@�{�qgh���MK�����r-�����V��7��\L���Xj��0�/�҆��N��pi�b�7��fŸ�iH�E"/c�fD��XwG%t2s��1k�3ꮡ%�WO��֦��}2ݲb����9����Go	4���,��%�j��'@w7�]ڏo���R��A�L����54m;��Dh:f�����uWn4Nw�>��P��:E�����.D�z��-����G����g�w�U�T��z��@)�K(�k�������F�e�=M�:{�����v����f���w�BZu�<�|�,U����9�J��XE,
@\���}��C����q���]��o��q��tLu�B��D�˻���i�����d�'�tä�3�g��Ӵ=0jg9q�w�4�c�Y���=˸4�N�K��':]�6��>^�H$��O��4~=/MY��~+���"ݿz�[~��6����:m��N�UoA^;�ĮL���RT �z�CJ�;R2�8��?����ޏ�oe������N��.�����=U�n�wwQ�gN���ʕ���M?J��ɚ� I�P��#m�at�G��N����o�Dڝ�ZUIװ�V=/IS$u�/Щ%�/n�Y�1��P��`���J��۲hԭ�BS 2=���bi��w��UZg�$Q�Es��i�t��.���c��i���S�ڶG^v�>�:��t�sE��.��M��2�E����d��0�cL64r/�W��Ŵ�y�����Z����5:�<&�+vU���X�4`H����9�[�;��]���y���zZ�b��dh&�[����f��[��X���h�ƞ<��z�9���?��hzӠ���g�����wq1z��zK��ŵ�>'L�KL�:4��x��E�%����𱶾�/Yz����ly�?K�`��?qT����K�q�N!�"�YY�2�����S��;/BM]����no#GG����vƋne���H	�(Ď�=^��k����ݻ�� �?rv�󟦫ָ��e۬W� M��v���g��#�<�i�������n1j� �^���i�oI4ZQqK6��+1�Qu�k	q�L&$����� G�������j&�D&c��P'{Hh��`�qO���Y����>�q��ӿ����>�c��xu/a:�N�o��e���Sb���?X��k.Ǧ��\J�VI&ŵ��ǚn�|gQ^��v��]�vi�jQ���]���!Z9"+�U�Ga��E7�)���:�S~5g�݃���ЙVw�,�4k"I�q�:,n�Z��X�<����7��];�����N��A틨�?�ܾ���r���4�m>�M��/R奵K�!4�K��!|���4�t���lX��S�mwE�R�R(�R;�Q���4�"D�ZbݱƤ����>����+�-n���m-/\�_��ڳ�
�%x;R�Q��Q<ii�y�&E>c��?�B������O���eu��������<ޚ~�������ˮK��'��`S�=)�����"�C��?���Mø+ŧ%H(ޒ?��M)�I�b<$J-���I��R������=��m���y��Z�v���]�����u�j��3}�������5�w�>{�ڎ����Om� �ud��l���>��lj��WK����8�*Y���\C��k��~��ٰ��}����qIfRT�>_��*��/�#�cp����K�)c�Tz��ѽOH���Zu��ͥFRQhU���.�Ȩ	|���Ha �O,#]n���߯t����`���v��]���SF�/d:[3�{m����:�R�p|���%y�Aĕ'%Ț�.����LM���[�55�*��ږLQ�-�VSB�j�B9��5�/qљ��ɛ/:�-ݧ|�W#��[��#Ї�5иx����Cq�p�@Z��c��$�?��Rv�B�3�+�4̌���;�����h��V^��ྋf�{y��D�x��>]t��F��>�/���ĐُʒD�e����9ia�<���#�S+w��J�we��5i~]㓵UӘd��{T���P��7��E�NM��Կ��Zvw�}��N?\���:�/�tn�i�1�b��[�&��b�=�c��Խ5�Y�NTe�KJ�H�$��K�c`����GmK��«"���甒,+ʞ��)���OR����ULX�$�}��Q��F��F��kv�g������Wi~�}�v�YҺ/S�1�w�}���z�z�N6V;���Uj2����Eedj����t����\a�#,�w <���������y'��#��G�q�&���?�����:5�o���Ƿ���5p�z�op4�t�϶�z�۴=���ʸ��8ʃ�u�dd���9\M�TUv��؈\��(Y��G$�f�U�Å'���CU��1�����}�� �?�G��F��n������X�gI��F4����n6˜�����C�z_�O,?�+��ҟ�X�)spj������nW� x��Y��~�c�馅�>=�h�<z���r6����6 ���}HG(� ��g22���{Q��[u�N��p;s���?H�k:g��z�W=������z��
�ݽ���5:=5�S+'N���d��+c$:ơf��V���G�>b;=�꼣)F����v]��xmҳI���#w/�q���znC/�A�}�U;��=O�D4�N��|S��wC�Y����Ƃ"ke�g� ��n�(�����T��� ��Z�bǚw����s�A=� �s��O��uz��F�ah�}}�'���^�K 4���b���� �g�q�����$�p#�,� \�����?
�C���fK&�m�j�M�� <9r�o������� !A���~y�?׿��f��1������� ��.�����u�j�M��XƦ���\ڛ<��?�a�����MA�5��=��~~�9�x� �T�F; ��4�j�������-����;Y�c�!@��rZ>�I��y!�7D��	��u�L�nW	�я�O�y<��Ǣϊku������������~t7���mo�]��M`��E�n4���n��ޫ��'�zC������陫��5jg��G]��6.��K&�#��b_��|.�zGOu�lӽ���+ц�JU��i�a�#  	�#�<�A�2J���όM��uo�zծS�`���Ob��V�	*$~ie��7D��sX��U�#����o��Hf�>��N��^�,�n���D���P��u'v��uK��;��6>5[��c�:�>Z[SIڨO*5MFkvB�|���6�Bޔ�'�h���iVZ���u=�ʿY�4�jU>�+�� 3"�>�&����/����'M�)�Y�oи��'���]����S�,å�e��r�5y�+1!ώmER���/��ԅ�Z�_jT܎C��;��/� 7)b2mՒG�qa�&��������_lt�C�ܗu�[^5�Jw��n��r��V��<1��sYd�c���:�z�Q����V|L�ONZ~^���i�weɎ����ah�UFb�%�TW��(�Gz��/��A0i�;B]���"����F �_G�r�e��;�oN���~���;�g���/F�|����2��拂	��/<?i�Ȇ�9ʴH��RKJvgy"F����,"�~�d�*�1�J�LlB��F��jN���5e<l�"Iu�,T���<���3�-���>'���`�_>BGM=�|�2SN.�6��ʲ�ߗ�ƠO!� RהT���w�!Qw�#�A>^jۜ
1��R �^x�<�Z��ÊrRIߋ�c�,cJ�R^Y�I���6�yE�C���,��;��|���2�Jb��-b��&��o)�ܛy�U��%|��{�,���Dc�5i��dt���#�9+L��X��AQH�8��l�.w����m����� �/׀foLd�������Y8~8��_ۙ�E)?��)%�_���+��2�.��7�_��E9]?!qw)xA /������1�i�o�7��5�c,��=L��������.����zcb2N�L_"�Y_!���锢g�ʍ�~l�x��µ����ͷb�Ĵ�g�\R������>Y��J�1���(�ER"���7 ��r^�yFn��!���1�Z3M������fb�u+V�;/��,Lչ� c$+&���6Y��"��wv1Ǧ5�j,'5��⻗b�35�9�5_'�2�)���X�a࢜Y��]�R��DB�KI�WZ��qD���� ۲� �W&j@ߒ�c�UW3�G�X"�p�㪱��izv*Im�`���"��f�l�+8&�k3rpV)���dgf�� �vcE/6[�vQ�g��/,�U��m#$�6Ey����9Z�LbMg�0�Fs�9��:N�}�&�E�#j ��Еc#��РE����Ĩ�u�w8�*����H @DLc����(SZʩ_>>X��ŤXl2�$���V3a�%�V����.\\�J_�]�IS%�J���F�0m�f0Bv��-9���ػ�V*%gE%��C�r��O��
� ]kC5���Wl`u��A�E&�`�2��c"~=����_1L_�u)�EAB��r� �G��`ޘ��K�<J�|}���/�VE�&pm�L�5uVFߎ�c� ���i5xʩEBnD���2,�*�n���2X��]����c�b$�l�TZ��h�1�%���U`�voL`�6Y�����,Wʿ�ԧ�I�Z��\"3�m���	�!��w��U�9�v��.�5V8r���z�]�iM�̱`�������'�v���(5KU>G0�쪞��Ǉ�1c�mE� g$.ʄΗKU"�;Rj_Dz������0���zN��ֵdL3�GqFJ������0M��Of1�~|�{bȽ�~���"�y�~Z���|o'�!X×yۆMjkT�,[fƔ��e_��*�,�,���
�ՌA�V��D㕎0�7��C�E��h��	 �mř���<�I�7G\�X�	c��JK�r�i����Պ�oʊ�,��R��K!
@��h$�cG�m�9a� Xq��c#ͲZ����bf�:�G�ɔ��ގ��(�5C)F1���a�
B>-�lg��DǤ�fD�
]�褊G&0�Jf_*�L1�#HK���5iG"5�۪si��}�,b"�8X#�E1�B*&�Z]����{M|�z錍i 7NyM@�8^�Z
��� �eUUV��FVn#qŌ�腚b���$�?�A���ʩ<��;p�b�F2AiӚ� ӵ��v�-S�<�c�f(>�Au]�ٌnBK�TM�&Ք"q+T�f�;ӛ77�U~�C ��^;��F��"M�,�sȉz�Iő���0�v�Y�^ c�
3dq��� +�%�ԅVr��2|�΅N;���1����<�,`��U�5,�oIO�P��2�p#dT'�c%<��.9V�d�,ȘD��
�eU0N*h�Pp.���������ZحN1�XPH�/�j�B��Zr%��'�T�3K'�I�ij�Kw�R�2&꛹��ߋs�r,cue.�d���CcCe��w3ɻq�@q��6	E�G׃i�"}�3nMkƵ�-wt�nb볣*�|(�e�Ő�?�+B~<�K6�uU����E,8���|Ls�X�SbfB�FPHV4���e�}��� �OϦ3�gZ�kiS5<�%�.V:+:J�� .��v]�&V؆�w!�61)%T�Cv�.2:�d�O����x��� m ��2��01Df��R�T�+�M�QqY�^F�a=���C�ٌ�9G�,�f/��I��C�%f�a��h�I��w %�2�<_hP�5�C���X��4�2g2���ȁ��b���#�Ɣ�K5����J���� %ܖ�;���fߏ$@����`�d��w���u�����f۪+N��W�I-��V2C͕�BEh��|�ƶ@1�>�]�(�.
���m�c*�*c�\�m��"�q׆߽E#H̃2��v;���<�W�EZ��#Gf<� Ty<��u"�K2���W���A��kL�R @�w�g��Jr@������c|q,�Wژl$�K֫T�W���r����W���ñ���C�SN�Y2J���C�*�]g����JѾx�c�ōV�c����J޶\le�4T.f9_�V���r�eWf0,��,�����x�fܕ�o�g�N��b�%? �V2l$�<2���^&@��OCǇ��㷒�_.�a���8̑�>���I�i?3d
�-j$+v���<��u�W�?�3	�* ����2����J�3���	� ��&
��zc��FvA�f�� %�7��|��`#��t��L�PX�	Θ�,X�q�m㬱����J����7�P��gf`��R�SɾN:-QyDT�@n���?�+��4��<@Y����Y�1�<�l��9>=��z^�@�A8��4׉��=�"�G}�ߐ9$R3u���,H'�%�����Ͱj"� (OՌF�Q$���#	�i;<�99`I�����O��c-}P���]C��X��~������R�6eI�?� 9+�>�0���?P�I�i�߸�g�Η�3��i&ȔY!uQ��e8�U }���C��ĝ����ቁ�8�� _��w��3Ϟh��	� ���`���D��l����|��5?�eT6�C�*��؅�N��T�G��㟷��Uv�(��7�?���g���V��6S)��g��
���عl7$�N�|z�k�\x��2�`O�� ��r�8oa�}s�����~���+Q�Jj��W�Sk �sG�<��B>?�$�Unҕ$�;��o�*x��}_a������V���Ƽ�|��߯o��퓵wе���/�c��-*��J�7U������+Q@c���� 0����#�z>��V�Q�7kp9D}� ����Oк�Λ\�}KP��'MNO)d��Y٥�|lQ�L�v�Y��8�UpO�Vĺ����=�~�v���s��<��x��e�:��Z3�O��#�yn8����/Y�����u}$��������iT�fe&Tu~��Ski��uV1��fWs��OV�uH֕=Yk��Q&4���%`���ā��-�t�V��rm?�lc*�F܄�� 7ן�y��������S�O��js�`�����DE�C��U�C�[6ŋ�d*0x�z���zK\����]�b}�����Ӑy̠��UՆغ ��W��@�x�\� �y��Fn7n����J�gVvg��GC��k��N��-���7Fi=0qG�n��,�=0y,r-��USQWϴ?#!��tn��MO���F}jv�������s�u�C,Uk�R�[O��b�0b1{V���cEص��t�����9�R)e�eT�c�����I9������݇�@wK�9��n]�힅�-?���H&�ؾ��i6�;ܯ��:���<��=2��m�Yg/������J���Ž�}սs��������]�sY�*4�#����e�Z�g��I�&�;1��)F��ST�[�Wt}�4���3gڊa�Q/f�4��j��	n���#ݧدܳI�<���o҃D�sOSk��;�;Õ��~��WK��;%��9�i��]gݾ����Om���8ִ���21b蟁'�lU׽�{@�>s}��-4)
M�u:��ie��!�EV�冐���iѸ�(P�'� �'�CI�����H,�ƌ�|���1��TE̓:@�{�Ա��?����]����i�c�~��s�}SPֽ��_T-��n/b�Rr��=�w�+3+U�k��������t��beY�8w����Ӥۭ��������0R�o���ꖤ3G�Ӛ(��*�kR� �,�UԈV=��u�uٶkU6�~�5-O�B��y��(�F�i'�K��m6	]"��*�h�_a{��F���v�?I{����R}Mފ��S�ո�>1+MKCԱ5�o}�˥�XӱQ/�����fu�}x�g��\�St�D���}��۩�AdI��Ha�,$n�XO!L��	�w�D���m^.�Ÿsk[U��$V���*�<6	�IdK5̒$���B9����}��2����v2=����z�R������=�t�e2{��db��^FNK6����F���8u���\y��>ӿ��\�u��.�T:5VU�WҦk�^9��O8��1%[�O<w;����h�V��"��vʑ�Qo����޼�O�����f���e�w��H�~����y��ߴ������`{C�~����u7O��u_��Xy�g�ײm�\{W"�|���ś�[˯�?�%�+�ge�:�Rg���:�?l��E�^�W��[���Z�f��Jǘ�b�s||ajR�[�i:2�թU�|t��$%��IH��3�I�7��(�T�vcۏg;{�]G��~�>麛������>��Oj���)�j��kI˶��e�Yr��q�QLnW�*�3��%}�_�V���O�/�nܫkn�+i�sM{5�y�����+�	�~;����ȹ��o�m����ek�j����Q^5�W�V��k5d�`2�A$@ȧ��<r#����6��N��~�=���L=o'�q��Q�'V�]�ֺ�矙����i�ĭS��\v"��oȥ.�3�36��5�[��Pe+XV�F�/b=���)'��%��UT[���%�t[;q'���yM�;�A�Ao�T c6���b=����o��=���ԣ�P�p:Ϫ��j�D�e�.�=;�� H�c�SG�o�gX�#N�1�.�W;?"�<k�� :o�Ņ��L4�Z-I|�$�]�r؎	�X�v�H��,�&V�,��D��wD�u?���P�%�.�
�j�1�F�璵XI�d��,�3�Q��K�<�+��+��ڳ;7�/����'y{-�?i����^tv_N�MT��]3#'T�'��Ɏ|�l}I_�y3���#���}z?�Zz�=N��3H�������#����R�'l�e�'1H�!N٫�I"Ef
񚞳|$Cи$��Q�ln}�ZΧ]��nԵZ�����3F�z����LN��$��_�Q��O�j]��}�{*�N��~~��}��v?W�:�O��c���>���"]_��<��	F>DJ^=J�h�Z覭-�,\�w]��:Ui�������ݴ�,Kw$i`��I��)�c�� �n�i0�N+i�FmFt��:Ƽx�Tk���Q�����a�CΎ����=�鈴�%�?������[�W_�z);f���X�_T�:��N��!�n�r�ˏau��طwTҫӵ,u4-)�-.>Eܱ
���bs�{S<��Y����P��/P�z
�kV�Z���%�/,aT+2��A
�1Չ#�/�F��>��߽��{�S�>�v�?��FKu�F������X���\�sT��n}��LU[����҇%z>��j�N�е�:���+7�ݐ�#���<SO ,��̚��Y ��F�W�B�����	�$ �̈;��r	�%w��^ͽ��O�u_j���ị��Y/S�f�oUv���+�۷�%����!|����5{W@�5a���^���H]�H��D�p�0�#� �!��97�J� ����	�x��9������;;��ܧ�mWZ�)���~��\�������׺�ሞ�ێ�H�Ng�6>�a��`"�c�)�
�td�,qF�w�xr?,I>�˱#���9fH��<�������G {$�v�1��F�qҚWI���� o�+�s3�g_�}�:����T�14,����1��=?Yk񪦑DL
���\)Y勶�.b[�������R�죉G%�
;��I�}Yd}[�YMR�3v�_�7=��}ܞ��'�yv����ݸ�t}�w����d�R븸�����*��GwN���/��g��f���%��|on�5m�G��0��yy
�v�O�e��{�����2��="�!����-<�!���&��?u��z#�zs�g�惇�]Ժ{� ���i��i{{��7/�)�5||{����
��)iQʛ�i�vZ��/����`Xx�������^9_�D ���Ь�J�9���'�����`y��G��YԺ����ڧQ����Z�Pk���5=O.�s\�ܗ-G�E�NjM Qg�د��>��˻ O����-K�.;�5��(�K�✊�@;2��������:�������2��h�F^A��7)r�-���)�w��r�f�vV��]� �_Dբ��c�^��ϴq#vp@���y�.���{�VO%�l�,�4������3��I�em�v�pkӬ��PG�T�q�~��2�]53�c�>��\�����C�t_S���GV�I�^V�y�b�y�1A��p>*�x��W���7YQi��K�	��qǯ�����z_�P���������ԝ���K�F���1�-�KI�]헧U��D����Ո��z�4m�GJw��I���۸0{G���g�Ƶ�=�HL�"��$v�>��޸�G�=���G}��>����Z�!��&g���h"N�a�ZV��^d���q>-,;�^�0M�3=�#�\���}py�.���2ӭw2
���s�G�l2����?��R��L�M�n��M7�t���M7J�]�A���u�Qk�����&��d��/�痒����rN��ek��.M{WԺ�NMjޥ4Zn�4 J��<q��*snĊ�YĤl�4��$鮫�X�F�iP�+��UZ�j7V�����v���7n�V! �*�J�!"���g���}���z�OZt�E닉�wA�I1��'RkQ][C�d,ƘY!Ъѿq�l��gB-h����@�䒜�_����V��Y9�J�H�3�m��Ͼu���V�}y�_T�;ݨ�wC�
��^��h�����p��һ5�h=?|��}kC�:��7*y�u
d�M�3q�FfV&nlg��3�)G%�n싲4�I�݌�5�ِ�cO������w�HLsF��6�Ŕ 9e�Nٳӭ����ak����V(uQ4^2%�Ed/ap�'j�v�t�v3�q�p��m���bߙ'��u��7��,�0N�t���6w�`�����>�lk=.���%���>V� �i��)3~#q-nO��sg�;�Ǯh�[@��9w6�E���хy�0���F�s 1Y
	-a��]9�}9�9:���=J�#��̥r4���$�y8�(k����x�`��j|n���v6�&��t+������A�����E��X]����t�h�M��4��ݟ�����;y��f��BݳW�����7���H�b�Ŀ��FZY��X�-2�XnY���&; �b��e#"BV�����C�x������qB3 �E �����`�0��{�/�v������+8�2,F�1�����t@|+""��h�u-4z֎Za��|s��TzcD��L���k5��2��011��gĹ!J}B��2���J+��L�Z�R���#�� ���!�' c%Vx�2�ǈ��+68��)E&A;�n,����2�2��p�pj
"�R��S`U�VU��P܍��O�0P�O�)�_{*Jx�!�G/  1�n#�y�X�v�a����(�uE���R�"���$�܏$���X��N�2rձ��w.�V6�FJ�b4�P;Ll�ʬ�VV��ͻ7�)���kN4�-o�/3LiFu�l�����P��*�5 zc ћ"���#�� +��t�^���]�dPIv���2�I���'TA%T�_�z������+����⛟La�柒��R~,Ti,&8��Sz5��<��"g��Չ�c#6�:5ׇY��#H�Ǚf�jlQd���@;��YW����9P�W�d��*����s�;~:W�H������cGe�^�"I1��RP(WjvfNqP)kBG=�X�:�PU�c��9q�7>`�pZ��,�J͑wE#t侘��n.Y1m��)� U64um�6�w�y��c����X��Ŀ��*c1�U���E� r��g@UKAf�~������9VX��͌Q$���H)�a]�´��x�x��Vӏ:�����(����G=�Ō%�]Ld�ғa�{	���!ak4	�<��qcq�\,���Y�Y��to1d Ԓ�%��F�$�b(��<\Q��?*g���ιli�m�0��)o�*P�$� ^L`�g��j��sͤ�.�K���X��t�ء݈c�����1x9QC)�"�p���I*��1}1�y'I�A�2#4I�����[��q�@T�*�bH�
�3c?�/�ƍ'F�*�r�B����w�˄�x�8�I5��������A�38���V�j��ͳ3�P3.D� h�˙�gi��x㌀&��Ɔ�Tݧ��\c(�
RCcjVGx��U�736�,�uj��"���Qۆ�c*���J��H���V��yɛy�uVĔ� k�� ��Æ�zck3J=�#4I~:��n�3(31R�WF^�� #+ �52#�m�R$+J�����TV��J���Ō(�H�Ll#�{�&R�3Z6�ͅ�i6��Uv<���*�P�dr��j��O�mG�J0C-򨼉f�YT�&��1�+��G �ӿ��o@�EeGb�*���U6�R�n}1�Lr�SF�Ǔ�3i�����2 �CB̛�3�.��1g75Jq�O9�P�2/�b@�3��5�ᙹ7-ٔ�� �h��ǌj'Vg�|���R�X<X���B�����Zc��2�&�!�]�m
$��AfV�����Av
� �;�㷞��>:�����sa/,yZ5�ri���'����dd�k�����*�9 ��:<�DW�E�ˈq��0�}�o��9<��mC'o'*�-(8b�<H?sv)�`���U�I���q�"4�;��u�"�j&\�M��b?{����7�0�&2�5��q�R[K�x�VK#��ll�(m�rp��mDgu��V��<��T4H�f̣�0�y��NL�Y��֒r����ay*�	+1�殶>%^G~,QA-��La?n-����Y������̉�7��څ��qc!|��d͑1�g����dcx�-�bD�F�hn�錗�����µ�ͦ���R�AEV���C�l\��U���=80j��]1����\P�� �"�'�T �59�jQ�D���'�‴��W@�,����žO�03����[C �#��,��d!LN%9?���[r�`���c�����P��(&��2!��NF�e<��R����t]_��T�É���-��ŷ����?�Lf'�ȵ?&xD�e	7S5���8dx�� {6�U�楌$Ҳ��~{�y0��Q�:��Y �"`l��o��0zdU�<`ʹHferȓU�Q�����PŕhK�c$S��M'F[HZkr��G7{d�^E�F���o���2*�b��wDk��,��7�z̮F+�9 ���*���taĐ�Ms�|zR�$���F�G��N��I'�$tU݅��ǳx���5�j�4ɿ�A�JYKС������X��g����⟚�c��~�t�Xy�sZ#��Y����M�d2&MZ����4V���Sjah�ύ�!���c�T�q\�\~t�c�%���&R1��GM�O`��݌�e����X0r0�Q!w��7U\^*6ߋ3��/ V0�����'e�K�%
�UU���B�l��(܀�5�>R�f��a�+n���U���cQ�cdE%�`�2�p���D˼�3��v��������8-�m��*Xʯ$L�;e㖓&8XG����J������T����U�%��Wc���Ulz-����X�q���+��
�G�A%<t���ԓJ�,ϓ����)�+������eJyl��yc+5n��W�A��yn�z�M�"�����O���WYykY.&-+y��qG/��B��<��ڬcl��<�1�h�
�>^F.�u'�^H\3�c#6�r%T6���ZZ�UL�)���� |�ر��"�b!�G99Sj��Π$��{LG�d�D�1*Ve�e��r�|h��C,�Ҹ�Y�թK��)ə���. ^-����ZLb��E�X�i�!��'̢�b�h��b7*�d	fa��$m�,���R�gb�hx��F���eD�U@`?���?�|�h�r:���$��h����^r���L�9� �iq�-��L��� ��%SJ����O�� �����"vϾIs� �~?�����jz�
�+<He�P��'$f5��P���R L�EA?>2]��v�J� #�?��?�G������Wh�=���9U#� �ϼ~�).��b�Ĵ�Qh�S��QR� �O��n}-�{&;48�G<�܏\��� n3��ux�/؁�������'K���^��H��	yi��d)���q��~�Ɏ�'�7�r33(�'�� ?��>����� �)伄��?�߾}g���~���4~��uJJ��S6�o��4�G��.���;Or�$�n�9�M�R���=�q�}�'�I�s���uk0��>Բ�~�?�{��]5S���Uj����6��ه�:���GG{eYe�����J��<���M�-�ތښR�4)��t����;���R?v������{iڛi�K���O�eT#7�� �7�� ��C����o�=ѝ��Ov�I�����k�[ӝW��}-�m���j4�tl��p�M�`��3)�?|��K��� wn�u����4�
.ڻb�QW�ti	y�Ո�Y�����n�m��V&�f��^*�@�O,�%HT$@�����a�y�:����s�����Oxzٟz��}5�GT췸�_O��zR9������?Pv���6��ƙ
QaE���IzgY��i����n�$v�\ӪD�T�5�(�X�KT՛�I ���U}0�j)궧5�oI���
;�i[��ada�Z�p�,q�U~���MY���I��*~�=����_�߰=q�||-9p���ҵ{��Uw�L��W�+��Ԏ��i���_=Ryb�{�Xږe�=�
��Lu���:GX�-�KPеX��mpCj-8�R#V8�j��b·�$.ѽy*A������ާQ��Sb�Rmr	g��\�ב�[AItk�a��V���)���x�O\׶g����}K�q�w����݄�n��޸鮚�r��|��Mg��s�j�6N��zU�hS�:���v�,�������a�;U�z��-��t�{L�G�Y���fm���M^}GZ1����1vi�trٷ0�uh{��}� օ�Zd�-M��sww�+ي�g6$5䂖��u�v��է��|�	x'��ݨ�>���<=�v'دb�+#U�=�� �k��ӵB�廡���/�:�#3/M�15�i�ȇ�]1_�J:�N���l��Tٶ7���m�ꚅ:cc
��i�׳��#��|��GRYc�c�Z���/U]��O��R�[��u�n�{�̑�g��� H�JT#�[�^��{;��;�O��]o����LN�{z�Ƿ޼�C�^>�=OOMcK�P�t��4����=�s�+�״�ec�d����>6���=5�ֶ�c�?W�r��Y�0�؍$&9�u�ya��:$R �@��V��v��M�oan&��۷��NX�d")�y�s.�e$v�Q�Le�F���i�]'7���5�-����̼���/w{����w�K�2�z��i8�oGh�С�j0c[��SW&���~��Í)z�����=��_��Ц+@��DJe̲,Hl��2!�?3:)\�����B�O�n��{xyh5��i
ז)�j��X�ie&w1�,*��j��?H��uޥ������֡܎��2�/�;��]���{'��y�d���ހ�/�jLN�9W5|Ij�3�R�<��SQ�-E�*Vy���&�ƫ�B6�Y�yo�w!���Id�cV��-BՉ"Y�jU�
c��y@u!�7�����)<fm��Xk��>6�u��폾�l8���b�z�?X���7V�uNcG�4:eWIi�R��9�0��㤕��'�� P�M��v>��&j:�����	^%##Wv��1'�2�5Y�i"Y2����kk���6��ܢ_��G�e3A ��id���ʽ��X��5�{{�^��?U��;��vO����%�l�g_�.����:˭���4�=�N�]O_�����cG6,�\����M�W�gM~�Վ�X{�S��P���j�׫<��bi$Gea,�����bi{���F��ܺN�!���R؂��'�Δ#�[6⮢:�D�����|ŻL��'>�M��轥�o����N���q:]��Ω��?�m=P�ZJ]c[�z[FI�z&6�ika�����W�}C�M����n��GC�q����0�S�g���,��ˆO?z�{K���G�M�Rݺ����d5�R�s��?"w�":���VE�bx°��5�g����0��=�d�=����{X�t��v��>���չ��j�&&7��c�Jա�c�>��� ��0�ot;�M�/�y��u��{Oq�$��߭2C^G��l��^���!�� @�L��D�����)쾗k3�p��z}�[0�ŉ�z��'� �^N5����S3f�����Xiݡ�bz��]��/k��_U��ퟷ�=�ӮA���ջ���W����/,{�P.G�ͳ��^��}����B��F�H��Ȓ�(�I��ƕ�(��VKA����n�������R���E�$*�+Q�[y�{�>�5���L�rJ.��� 5�i=�S��_[�n��u�������&���d�����t�j������3R�����	��)�i�e�+kR����K�<�N�c?{0��BWd���0�f[Vۥd]!#�l Z��(|}�bX�{|]�R�B
�*�f?���^�;��N����_���ӓ���:7G�]u�|�<�{�4�uH���m�SA��p^����M��}Z��>�"�'��G2B�Dh��W�O��E*��H<�GB�v���b��7 ~�AiP�/^���[�8K���:���Խ���V��k��Z� �G���z�^Ac������"�T�NW:.������ȑ�D���y'�Q�V!��$��>�V< ?�>�"�C³� ���>� o���O=2�u�Zv��=a�ڟ�\��}��5����t��u�tv���}7L�ŗ��ӝ<I>��k��/�r��  ^*賚�ݘ2E��+�~�/�`�!X�~��9G-�i��,��`�/�K\c�c� .���t�=��8�d5�SB�}��]��L<r!|<^��ɖ��z��sGQ�˝���*=^MK�\"z����v��?��̀�!?HDf�� ��[֦ͪxm'�u�A�+w���?I� �R/p#��k;�ۮ�jz��op��c�����g�=��z��SX�r��_ڊ�y-��4�T�u���]&*O'Q�d��j�<��(8B��ob��V@xϠ{�~y��˓�T�w�~[������	 �'�d�x ��5��>�޿���];���״i��C� O4K_6�G�>"�rz��_�u`���L��ci�_ն{�.:I$�N�C���E�g����e���^�^���%��?~?A� <Ջ�qp�Tp<'u�HP�0���� 稅�^Kz��?��p}<��c-�F�t"�Ŝ�w,���8�@n[� �}����F?e��Ϡ9� /ן����r�����l�"�/��6d���K�
1}�Cd<�������b���{�S��8��3��s�������qt�=r��?I�r!KAۘ"B\�>��6w� �����a�KP��z������ �|�[Ƣh���#�� �������8:��<D�a�aab�^�A��R��w�����'��f�� W4�<���y�#����� /�Y�֬')�X݉U�=�R=�� ����=k��1q�^�ԫ�eaVx��FI�X�O�ڦ\$^�!���	�P�a����R��(i�A���̢Fn>�r@�8���dZn�F�_7�F�Ğ�C2�x��'�G ���;s�N���=z��=�_#I�\}K�u�k#E�I��ŷW���	i�3��R���r3�<X�q�]7�m���ëT�5���N�X�+,�$}�PĂQQ����k�[I��֡�aU���r�E,�㳵G�%W�~�ߏ��?B������r����뮒�m���\�q{_�>���P������v�04������'��5gQ:U1����D��B�F�]���}���ZɛN�Q*4�E�1��Vk�%�2�.#&G�e�(�$f��:Vz�Srm}�~�ٴV-J�����kG2�������ZC��A���X�r�Ǽ�g�ӻ�K��x5~����>����/���W�:���;J��B��L��G������:�n�����E5+��9��[{^�jm��w���ĳX���HYf���I��<�]��E�$�p��A��
-6�ˈ�]���޾�:�֩[qU��zu� �������q��s��IT,p�倪F*�ο�H�Zi�w��O�eC?K������'M`��';N�-SR�5�!T�U��y+]�OW]�𷽴�l�[��Փ��p�;���d������Bp~�A���v��&���)Z��Yd�=����J��0�yIe^@�
�h�+U��Z��P��5>��-\��C��Ͳ�'��������v�����b��0�Ƙ�b�7;���������д:b��IHD�bĳ��yg�W,�Hĳ�O�i�����׫\ֵ�-f����BF��H�@���*"�(
v+�`���;���;'��۹ݿ����^�[e��ևKh��U���/#���u,�yɀ�љ!%uȼ�����Ԯ�����:�(�kC<֨��'2�$S�g�#�^�"�u�>�H��tK���=\�W��Ūv�
7^�0^=�+"S��RIx�[�<��������+M����ۅ����7ztMo�N����5�/�}��/Ѹ?�bՑt�u��M7�31p��Y���c�d��t�G�xt��G�O���ߧ[ܚDrG$uuV5l��(!�΂���JKJd�1���W�_�n�tʵ]Gg^����H��gM�V���}� 10�D6j����RB��ܒG�s�:O�[H������Ti��h��'Jb����H��i�r����+�,����S�=�Z�t���Z["��T쿵kr��!p+�3��Q��9[�=)������۝H�m�Udh��a4�\7j<����i={&ZÞY�_C1�.|%�������I��Ɵ�����l߉�
mi���
3$�����=Y�j�f��9��7_E$�º8>������^�{pCj��j���:�����"GR>̬A�r]g1�Y��OR�����ҷ��bբ�� `�O�e>Y�ƌ�-7�&�,�*��.<iv�ܰ4�0�U��IV*a�'4�2�'0[�3~q���T�y0��d���8��\U�Td6N=�#5^S����<�ɛ�e���q��2�K١I��Q.OH�x��X�&\~Q�_�I~�V�/�Xư�YK#
Qc�e^P�w$I�#vj�f �
��8��R�h$/3"�X��Q9�2�7�&�I�n@R���UCj��YFu7>b�h�E;
�� �f$��V0������Z����L���Qa���$���ld��C�EW6żj��@��\�d�P��M��/�2U��Ye
�c��sǼ�D��d�uDv�|A�g`�U�0����K<��',x'�y�:M+$���N܂!Ys��5��9cw�ky��/����Y�9d��|й,T����.0T	G�U�2h��M�E�2�%,�~)N.�0��y��9��A/*�?5\j����\|��� �c��D,��a(yy'9����<[�K+��Lb�5Tm�|����g��!�Pؕ�)J���ʔe
���c|����W��ֹ�V�4�f��5`��Vu-60�Uyc�,qP<[}�	=h%m�"P�É(F� ��O�J��_�)Ld�L� oplM*#*#)���l�!�I��C6k+
2y!91qQ=�j�{6�K7cU����٘�7�q@'-9��8!m�n<!�1����9�i��7�z,�%�X�=Y�ж��wFr��1�O�Ȋ
#�r�V��C\�6?�����U 0em��}1��X��&��_���D9y�:��>YX(�Kl�Hu�G��|���1���r�y4/��v�~�� s݁c*)��'G���~=���Wʽ���y��'e?,	 ����~,��Wdo(q��Qh��ӕ1鸊�׊��%�&꼷c�2�YYD,|���K5� ��g��*��U�m��ܦR��3*R�����n�e��S� 
��Acid��J�'$r
�E+,6R�����~�7(��kb�L�􈥱K��d�ɺ����LTc)��fw�(���HV~Way-?")@�����Ӡ\�(fA@ۂ��2S�Ҵu��]�`+��g(�Z�����%ߏ�S���t�d�E�V,L�j�I�j�-�|x���B�#�ȧ�1g,[T���'��Yj7��oO���e	��n~�1�����ҹ���V\�Q��#L"�b��x����KMR��5W��Ȓ�����գE� �F�O��>*LaѸ������s'y=د.M3ρ(Ae*�Pi�rl�T��l}��\%�Wf�y+�}���������X��79�T�F@�t*����i"ɼc&4����F5&��n���e�&�c|�Z�\��ɫ���$��/;��P�}x�9M�f1)�|���m�ȟ䡢�QX�s��*� mÛ��'����e�Q�Y��ζ�R(�3r��*� �B1�7�c���v�Φ51�|]���ro�>4ri�`�{1�
�̔�TR�J'���YJ�%�*3n��%�}~��X����� �xM��g�
wDo�B�O_�bQh��Tg)���wc�İV�!J�,dU�\�
�t-j!R�e�ش��,p�-��2��aI�KM�.Y�ڙ�o��� u>H�Q~��k�ك1�����e�='E��1�T�� LAUq0X	�yf00�6���)��g9��h��9��r�PO�ٌ(��B+*C�e���`�raT@I��
�e>=�l��5Q�r���7��1'�e����!P�� ��1c."@    ��@�  �ߙ� ���Lf ��&m;<yџ|8�5leC�sGTw����W� c&%$�EO��xǛ��W_(��1�eg��N>�]�2�֓��ŋd5����IF�g��G4fr'��T�������i�9^G%G5
�בM��@�9O�OLd��ư����ݘϒ~?�y�rX���$�B��(V�v2%��$�q���3�vt�3{�9��5m�PI!O݌�uu�6��:S�ڴ|v���eD,�W�Ň����x�Y�q�=���ɴ��]I��#؟��Ա�Z�#q����cYRK��*+<�S�y [���������e���Y���Dxȫ9˻��+8!,��1�^�ZH2דUo��R�h�v��ڋV2b�ERy8V<���JY�fȢ�e��S*����S��א��Bǋ���Tgu"�&��xH#���ѿ��Y���8� qs�Ō�||�id����[�w��g��t�(�*�\�����-��O-�W���e|$.�����2�n���� 	��iT�p�Zf#̢�T4jН��J�+� 
���1�ycH�,�GD��SX���� ��Tܱc�~G���Q%D���	 "��ą�#"�����{�M���A,c�K���z�@��n� ќX��r����+1�RBoIMD�,"�e���鍊��w��,��;q;��?"�gɍVe���ǤY��t'��\�4,����?,�"�m���PK&+Ή""���P�~w��l��
y4ϽV��<A�Ec�S�g��JD�,�>�QQ쁇&0�^2JRE6G'&��6�L�%��4^j���U\Lc�@l��BD�"/T��7��36$Qټ���� ,�M�qR���9�a�]+��˻�8�T�T�I���G�Rz��N�1��ӱ0p��b��sB�qe�lv���*��������6)�VD%H�(�59G��� ���W����Ry������dt�	�U�#���ˬ�oR�;F՛�6�������:�K���jyZ�0��gYKD\��%f)�ձf:6�N�'2G�]f!W��uf~A!H���޼��{�Jݯ���E1�q'�y����Y	�v}6������܄��'3yc����F�I�����;��,���?#�G�>� �9�`k��1����?�����G#_3xھ&N����� Q���9_N�f��� Ʃ� )@ֿ࿑&��(�Ν�麨:bjKWR�D��IK�;RR;VO��xo@��u ]Z��$�'�CH�{������� ד��4Vxk�֧���W�B��pru�?;��!��gi�����O�;��fIm��)�4�4��v=����*O$q�0%}�	|�p��DW�ي�^��$+G�������t3���u��w'�}���^��k����-KG�а��M{�zߨ0/���#f���8=S\�l�,�e���*=���0�� r�]Kv嫤�ͨ^י�ymB�p@�D�-�B�H�&Bݸ��Z�� ��fh�?_FXD��:AH���E�{e�[J��8���%%0����t`=��zF��|;m�����@�Y9��9��:և��T��	���{7����v���S6}Q����0_P˃�����U4o��:�z��{��Ey4=�Z�js�%�P�Y+U�$�Q�I�ZӐ��[ZڽA�֥Cwn����+�m.�r�����~��NX!����R�#[�6�L�N��"4���~��m>�����������o�s�k�]��z}�M���{:����-�c�~sq5$����p�xc��b��[�u��'�\ޚ.ߗG��<��Z�Y$�H�a�?�*2��X&e�h�nՐ�!���eЪ���ku�Wu�Ɵ56��?��i%�	�9�s,sČ{eg&De����=��S�{��޷��q�&1{eў�;��fk>���u�~��<�����o�S�6��rښ�.?J`�g�b�]�` �zW��ҏ�Z��C�7+����F�i����#T�^�ǖ-O� �J8��S�$�8�'B ����\7-�ӣѭb��QN��Kr�9j9����&�j����!����4���k���>����߷C���`��wݍ+X������w�<OU��ƧJ�/V�6��t�V})ռjf�����m���;�.��(�t64��۬���������kE$v'�dy�bf(�u��[�ީS��S�n=���Ef�Cc�Y��f���J��Iaq�a�@�Y��LN���w��=���W�foP_�5��'��:�Ժ�U����gW	:w��f��kC͕�`Ӽ���u.��W4�fW��ԟo�9E��w�X�Dn�;�,J��(oc��E�o�՟C��ݗz���m���#��� ���G�ݾ��}_���E��,�E;�m��u�;��{S�Κ� P�V���yz�p�k�'�yV(r�S/"n�8Y6:v<TH�ӭ���L���.�n�4�j%Ȓ�NխP	&�k$LcG�
����I,�Lm�zU�~0�i���7��IV�j�J�,2M+ٰLq����w�R�<��1Ƒ���K���/M�w�_ҫ�� s����?;��=��gG`b�ehk���C:�����cf�:n��S?%R�ն+RU6���u�#�z���j{;w��bZ"�;4�����M^���D�)x$E��*n�J�;�zC�ݻ3\����9�?1-;u�
��X�$�(LM,H�sD�/�@���[�� POj��[ӽ�����R��ԉ�Z�Z?\���W��kn�ԻT��z��Fwqsw6G���=d� �O�Z~�����.�ӡg1�h� �N�.����.I"��
?��o���h1N�$��[&0�G?,�B���=�(� 3n:���I��iߪ���]w�X���n��d;&0:WH�����wEѲu�̤����к��#�
p�:�gg�&8�z����$�_��4�Z��nl]���v��c�<��c��*��Yx튼*�[3�t'P����Һ�}-#�:֣�N�>�ר�]��i-�;Q1f2�)��.ݫ��������?L��~��=��׉��Z�����ҵ��KOP�5'�&n���Rv�Á����6H��t���]ꍺ�?�4`��Ctۯ�ޭb�U� �$IѽfX�P�'�22G�Xל���L�Y�e��[�@�oR�j�ɬW3P��	�ڻ!x�B�|L��*K�3tO��~���?m�4�i6]���&����^���Ɇ6���eO\Yj�D�?�ɑH�+.*�_T>�zQ�ϯ�ln]U���U���;��C$�Y�^'mL�byt�J9��� MҢ۴�m��p�5;Q��8)�WKk�y+uX����9�g��;��MW�������}{����J�+>��t�CU�U[���}'�LM5�(�e���h�>���:��_G��ZV��D�+��V��ym���v샟%ɋ��Q6�:��j5Y�T����Zω,�%�X*�/��Dob�4��ffw�]��/�߆�.�wG�tމ���Q����S�u��Ϩ�=	�^-s�C(d�@��[c��%ђg���UR�5�8Ԗ��E��}��	f0	�겯2���d7�.h��p�J�s7��?�b}wFYO�vYî�wڇ���uŻuԩ�ۺzfG���ӵ�I��٬�\c����9�1t��)�k�L��mX��(>F�l��ly�ܿ\X��K`���+ܧ��:�#����N9y�fh���H�p����ݪȣ�h㻏�� ��?j��R.��;��ί���5w۹���	�O���'�.�ӓu||hD�6��KI�Xx�'Ut5-ZeXcg2rW�fn�I?`H� l�i�8r/��� /�����󹽎�=��(�>��N�iy:Vu���#�p}K��n��u�/M�^���AʶWm�?;�1�zE(1%�}/Lzd��2�x$U�c��l�VB�tY[�2+FH2H�6�u
�H̼�zY�^�dr������K�	���������r}�k] z�4��S�K+F����9W���W��<D���(1߃R� d��)/k:ޜ>Ek����E��w�2p
2�k2��E��}S��]�%�ު|71�������q���*x畺oqtk�f��E�>���a�Z�]a���]��-1�g;8�o\`�R��Qq�*D��0}|ͫ�0�a\Ƽ4����
�آ��I��?n������I���n>� ~X� ����FjW\u�P��Sj=i�G�uwV���z��2o�j��!T�@%Ȇ4�B*�e9��c������?�۟|�I�8�=���|s�� � �<k桭HT�p�\�CO�$(�;� ;o���~��S�r�?�������Q��FZ3�/�Z2Q���8nU�ߏ=����  �� ϯׅ��Π0�q����� �~����'�G'�i�>���NK1�(e�8`VX��ܝ��m�ޭ����%�@�8��?~����P�_�v�$���� ���='Ihٹ9�0�ƍ0�?}�#̒4�样.�����]�n²�q�>��G�?Ny���e��ڼ0�� ��� ^3�i8��9�r�qS33>�cRSn$���O�>��?>6 l|��=6��+z��z�������0�m��~��?�	�� LL����{/��KtW�k���"F�Gԯ�3�h�8T;�I<v�ՕwN䮭,Z�q���<H@�$~y�����˓��L�$���$���|�>�Y���L������U.�������u��VQw7N���-WK�N�uv~�n��0u-#5��'��y:Um���n(L����N�տ�ܯ_O�F�U�DZAʙZd�\�a-�׊� ��V���؆�ӝ�C}�EJ#���"�A�3�{`�v�'~"+2�����x=��?���4��s�ŵβ�z����}�u}zc�]��^����n��t5ջq՚�MzwO����WG��~>.v��c�Ӗ��~���4Ɏ���i����$w���s>�,dUԤP%����^B����vuqϢ������E��j����#�#*�ԍ��X$9 7F��w��O�M/�}��E헯��uV���b��u.Wm�u��qz�q��_��'^��35�7
�3Y�>���	��POM,|_o;q�w6č�R_a^��ε`i~N/�����JƱ����!}l���R��lTM~�[��$���2�/^y!��WH`dh�&v�ńO3���=�����@������{���O���z��^�·Yg����5u��S�R���0��&���Ŗ����!b~:+֍#�[k^�z�[�>ߥ�[Y��J�b�,B?5aE{��Vz�$��Th� f�u�z�Gw>��t%�T���i64�=��T�$�Q�"ILt��-h���BG9���{i�K��1ғ���{��^���ot�=[�O�ϵغ��p��R�����ة���:.�|�+���i�2g���I���ww'L�՞]�g[A�y㋾����9J��j��a��)�K�z��-��:�j׶)m�]�
n
���I$�W�F�v0��V�#BM��M��K�݇�:z�F��lM]��=}'�_�}o�܁�	� mZ�N�7++P֣�-,R�G��qg�-�n�|e�����2��V��-ZӨ��#�Ԏ��"-Xy|��#o7-��� E�:v]K���3��)��;��F{k3]l� �C G �m��Kѽ����t��q��ُx�Ӧ�K��9�z���=<j�T��<�ፋ,�Fu���Irբ���΅�t7�Cy�]ѵ��՝�n�B�[�ɪD$�F����Md��ц�$��F��V s���e�=��]���e6��z�	SJo]J�qy~hT���B�J���,l���nz�{��%�Y��{�����uWtΛ��i���%��aK\��ӺoL�Ma!�~MY-0��P���T��Nv=]W\��n�:��(��ű�
+�$�$��Y
7��<�j=m����m�� ����X���"��I��l���0��q����+�$��߹�￵�S��7�?�������M���U����qp����m�k�v��.��LOl2-�.cd�՘(�
�[:��A�Vޟn̢@|�SP��(�|�"We�Ohl�)*��ڑ��'Ez?��-O��CM�F�!�-:�8C�,��������ǰ�<�ү��L�~�����i�����{��v����^���WD�F���5~����M�SW�-L��u�G�lF����cض���u��=.���^���&9&j"�Œ�e��^��/ˀ�^/����^�n=�'K5H5�j6c�J0��j�r����bU���7�b�X@�K9a2�ں��ُ6�S�=e�Y�3TIu�O��F����Ti��ޭ������FyX�dT��'R:�v�,пS{m�ğ���v�9�oS�I,T#��q-n�� f}�N���^�}KM���%��P�`��@9"�Ǎ+������Vaփ���_jI8׀��8��V��v�J����	��#�98}�������i
dn�֜�)��$"���p����T	��X����@���Si��w-��<����M*}1�\C���e�R����`�{��	�b�%�JQ�V�����vx��s�rx�.�����O9��Ʈ#g
���?\��<���e�#J�Q���8+�?����mtyE�pi�������!��B��l��w��I,a!Oޡ��U�|��I��(Y���?��������lq�θ�x®�8��l�ԉ`���}Xr�.P�2KIq��Ι�F��N�U@�Yd��I4�M���S�\&౅�1Y�=�Ruɢ�:�|$�Yh���*^-��!@+�g��y�U����Q9e60  \̓P�+�ٗe"6�7I�3N;D�ΈTHs�A�J���<������Vi�͟�k0�����`���0;�c��K��rv�	�K宼� #�-'�L�S��.9�C+.���{�ZA�8��8M2j����V�R*�Sr����	"�djEWr�z��L���3�ę*V�	Yȟ��G�1,g�&��%�jTs�8Х9��Gf�� j1$�c�e��ԭJvs�(n�G���� ;��s�cs,z��-J �֙A&����#e��X0�&i0C/ 1�se>JP�n�29uR��\u��?Q�w�慆��1�y*���+kD\�l_3ۛN��Ŝ"-Y��*��`�.g����$Q?d�';�P`S(�� ��j�zc��J����l��7㴲Jbx.&�VW��Y@%�rHH��0�&�ݿ����4Q9��+y��*&�=8����ı���1�f�ݍ���2�W������u~"{�+x�U��c?(�+�.�w�,_$���1�~�J���S��B�12���-��>�oM�I��ʟ���f�g� O�0-�޳��)��U#�OW����Ra^$Ki�
���zc
����Q�d;�^��p*�C^�$��3,7vر�pc@%lJ���75h�Я'�0)ɷR|��|�nX�{�T�X���,)4���p�zrR����	�t#�2S`��m�vZ�51�nr$���Q��*ǓU�П�� ,bGcV�S)�4h�:J�{N��� j۠?��˲n�	׋���ҿ�d����,KD
���z*���c$&%x"&;dC�&�lJ҅h� �yx�+ ��cJq3�ǔړ��E��L[ �~W�[|L��|�I#qŌW��T>`7�����L�����nS�@o�N���n-<���-���eN��Ḵ�z�'e񪅐3
Yv(Ǽ�fc�/!��|��UtF���/�;��@,�1�xmY�x���(�����ƽ����E
A�� Bo�������ZI�!G���Uy�y1%>�Q?�OLd��?��� ��D�F��v�%t����B�s]�2p�{e"�e�y��5\U��<�93�~�f~��ٌx(N.<�/ȭ�S�*���G��6���łWo�c�e2Y��Y��U(�J��Qy'��*7#�'�%��+;�:�P�ʼ���3>=��He��F;1���-�Q�e�Mg�mWI?���O=8�Fm�K4Ϧ0�.^Z0sR��lgt��B�4�!�D���O��1���O:�c�-ߔJ"Ҝ%a���~0!�䉺�័c$н&�f���
�OZ=(�`f��V�"B�c��"��.�L��,Ũ��S���fG7p���0�R�(K:�*�j+[�29e�)2����Ó�~g5����-%���˾6�J"IԉѦ����AF�oEsQ�B��F���Vj�rl����i�Zfj��I��ܕ%9�1�xN�%Ƞ���V�b<�X��t	�9*����ac9��lz7$y�"2L�[j���U�+���,`�>���e��� 3a�P�1�m�����N�r�W{RA��#�\&1�_�l;,����2w�M��U���r����x���fH�y���Dlc���P��)���-Y��;K)�%O�c�QjȠ���)��2��E��8c��L�v53�kK=5f�f�I~'�3�ԭ+�g^N���-��N�$Uy�2�vG^.G�/.e�����s�ka&Fa��2B��B��I1V�}8ߐe!P�Le���Ph߾Q����|t��>b����-B� ��@�X�����"�(.�̄���f��k���9��;�	n@X�t�����eP�U�c1I�K�|o��5*j& ��s���I�qE�d���"3+䩻>5��B4!�`��L�3@��+S9H�UFxN0rd؍�d-��d�b���(�G��	�1��ɥ
>-1��2������!te	�	z�+��E*ޘȥsc���dedu*��;�-������K�lH��N�Zd2�.;�������:�5�W|:���@c��_+��C���gN��d@�4fm��7���pX�����ߑ�ҹ��$�b�`vI�;��W��Ō���Ғ�ِ�>� �L��P��A��4u�E27�ȏ�)
χk�ޓ��!.��H� ��1錗��!|<�)�a�|���5L��	(�S"�n;wf�X�X���i5Ǩ�f�ė�O����NI�� ]���cI=���L6���[w�l�M��&�*m=����02*�L�����'�)�J���i�+�d!�P�ۅ5@]�1��͌h7�6#!h��p���2E,��K!J�e,a�*�|B��:P-�<(����l�0�4�W
��~*��ʊ4m�%4|O�ȽcK���u�y�ǃ)�_�c�;��3���|���'/A��֍��g��}��.��ka�f���m��U����4Xe�dj�����"�R6���X�9�����S�-�#���pS�w��LQyXك�� ��#�?��s� ���st
j5ӴM:�k�r���]+SDʆ����{�W�6�&�F��e��_E�"��۶l�����ǔFQ�~���9<�{�O��jZ��fX~Y����8^��I� �n �@����J�]3R�������_Ů^���"
U��u�iӕ�$��ި��MN8u��_�*�P? J>П�����ϼ����:F�5XZ��?�1�q��!~� q�=�d{a��K�S�v�E�N����t=�u���2�_����2ņ��:����H?��O�ċ:��z�s�V�Gakh�dR��f��x�N�%�U%c��o�7kVZ�z�]�g��ұւ2�'y�#�O+����Q�y�';C�O�p���/���V�����^�ky�G��p�S�����MG�}�k�FF�ԝ��קK	�cC+Q�Pɚ6f)��\����Jz}�*��ɬ��í�>K���u�b6�G�X�j񭘕}+(|®t���v���^��H���,6㑿w�z�;&0G�mwU���ú#���.��� �{��N�wW��OV�c���n�մN��Ś=Hz�3R�n��m[��@�g�~y/��G$JZ�3٢��o���U�h�a�[�M�6��ji� ��b=0ɧD��U�ogE���Y�5�v�y��K���}N��MCUؚ�س��R�j�i�X��Qycy�ѵ�W�^_h��;q�$s(
�<���h=��l��'�k�n�`w�^�z+�:���'��5߮��-SA�4oo~ݧ�MF���Z��ԽN�}3���Բ�	,�����>�)�=ú�m�6
ǭO�-�t�k	I"���/J���%���^)%�*w�\��4:�{Rۿ����?i�\�%�c����$���rĉ�d���B���/}����dv�� �g�=�vK�O����1qu�o�8�Q��Eԝo��ڔo��T����������f��3�-xβΏ��n���η�=�?|p߽�����-�Ϥi��W���Փm���'gS�\�`�:�ڗN�ux��ߝy��F{sZcڟ3r����>Z�˪*�â���bź�羮����Ե�/���{��^��Auv�O�����>^��lmSM6�ϕ�3@lf�/>y�y3Q&�� ����vѫ��n�[w���T�XX����D"�nb�j�E�,S�#p�ʅ�+��dߟz�͙�鵷.��\�2H��O7|�]����E�2�,3�o!�·����Κ�?�?��7�z�g���moӝ��߸~�[����zv�~���zsI�qt�����Y4lI[(�2��%�S����í�N���O�f+�P��!{P<IM�i���� C�!�B���o�}�ֽF���zmV݆jIrk|Q�G6DAP,-�Y]�c3W�"��O����~����=s������=g����뾯��@hC�����H�z¦���z���J��La����g��
��IF�c[�����u1��z������&�]����ei:�7o'>�?���������߷z�q2�lS�� e�*��
��F��YdB�# �3o|u�W����{��j=�{>��w����v5��t|�����еM!r��j:�g��AΡJ��A2�q̣�},��Ҏ��hX�;�m�4��]��&��<r+�v]�i*I�1Ⱂ��a�R���U�����]˳w2Mf�������m֑B�eYd�H剤+b!��<����{�������b{U�[����}E;��])��']u��n����$�:���"�:..\����s�1�m�:O��L�v����Fk[����ٯZU�-�,pS�~Zw����*� �>�!��W�f��SԿ�}ţ��C�u�ԥ��<4������hb�׎Uo~W� �/}��!{y�T{o�B{��K���#��i�,~�\\|^��s����=1��8~Y�^uᶟ�A�#Y����� H��շ��j�锣��O�ԉ�s^A�3=�"YU�y��HTspt_���)��j6���n_��-jV��G4^H��_H�ЇX�0P�H܆̃�;����Q�ƙ����u~�����_u��~�::��V��Qi�1�|mD���i�gJPX�C:v�m����a�u]�Ս�������^8kX�:�46YF�!���VXG(��]Pi���� �/x�Z7K5y����{5t�&I�U�l<!�%C��謥I�^Hx^di_[���ϫ���dvg��;�=�莶�1��=�{`�?�:T�f2S��[dc`�ˎ���)2��O��|BK�OL�j�.��n�M'n�|#�ZUR��54�"��^|W�F��'j���ԪS��mթKP��Ti��1���ǚY���=*�D��)e��떓�ǥ�D�;�}��p�+�z~���=1�����_�u��Z�_H��в1"�L�D� 	�y����7�K�_�5-A#�.�w���0��i	�!"�G�>�FU �+it�äS�?Oo�Z��!�UB��xX�V+�q�'gr�,u�ާ�jZ�k����>��C����J�������O�c�R/���� k5�b��c���8���r�)6rk�p�Jr��ҳp���s�:�� =y� �n "^���GiȩɧZIfJ�9�V^�<r)�ɕ�^�}����p���z��?������]sП�����ך6���~�;�$]B9Z.�:zm���3��nT�m"R�c��%�
ݖ�KSڊ\�:�׻�{x +r��_�ف�s�+��##>�8��=�`�s��/�nG�ң�=�׺O_�Ϯi�Sܝf�p�k�!��'G�3`��w��^0k4��1Âѯ{�n��z~�5��R"�5vWq�9�K�Q��ا�J�#�r���FH�=�H��
O�}���>�<gY����ݶ��ct�]7ObtG,N�t�����iRŖ�n���N��=2��cJ3��.��+؍Vj���q�{�>e�]�
JJ;��og-�%+�`e�Y^�py=ǿ��I׎xଠ��x�:w���{}��W^�Q�n��{ێ��>����CO�mk����cκ'gz(�:�U�Q�pt�j�����t֒�;)��4�R�u]ź|H� ��y����Is��	#�7 \'���K$ơ}�@NTV�� 9�pA#�a��������{q�]?W�?bK�~��Q�S��ȿ�[_�~�!/�YEN��(h؋4U�E �{v�z��e�����(�~��\����>���ujDU�	_��7���nx��5W+*x��c�N�Mf�Tp�$?��Q�v��o^��y�	8� .}����8u<_]�� ����]CS9/�\S0�Jxј/���̒H�~��[LEf"^C@��߯����?�S��zy#���.�:h�*���9LB��t
G��ݐ����-�6�ArŚA��>����z�?�ʘ���k��� w����9n���l�>&�J��I:l�Go��������+�H�^e2��w${�� <�x����=x���� �d\^��rt�,��a`��~�UVݘ�<m�!d�}�ݟ���m&��;�}�$���w�2�����>����^�{����F���5��i[�ьެB%�Wx�?����	�g��ڭ2T��  0f�?��_�?�[R�SF��_!��_������z���\�i=5����_�ܽ7'#ڦzc������+3��/.��ڳ�x��jj]��N�?S��}����=}���H�$mb�uY���I� �����ϯ�7���i��p=w�Y����v��WH��.������h!�wC�Աg���{��j)�ӻ���p4����j��z�<Y�le��ӪW�w�K���U��čoN���X7k�T��hO'��1&�Ի1MkIi��j�i���(�,7/��g�,��������'a����{{����J��F�ct̏q���wz'T�{ߕ���oR`h�--
:�b��P��㛩�Xf�P��:��E��.���^��
���N4mgfA�[��/Z��]��^^(g�nʹKI�I�z��h�Hf{��.{WiM����F�ƙ0��$0G�k&�pA:��4�B<��c��]`h|��za~���~Go{'�?s}��v��u�Ǻ���Ի��_�c���ڗ�.��M?+�Z>j�#�1��㍍E�w�����U��S�u;umz�w��sKӫ׍����4��gM�	w�zr}��
��r�7�*#�R�։�S�#��k��icnP�-�,An��wU�G*r ������ì2�K��{3�:kٟD�b��C��_ھ��ǵn�� F�,�?/���y��:S�p�ϧt��_BŽ�H#���E����gۭ����PhA�E��̴��%���Q�Z�3Fz��Y���E2����T��y��6�U�ǧ�vŵ-7�R�si�5�"*��2ي�b���b���$}�B2϶�{�)��~��=!�^�dv3�о���v��w�������f�"Z*C�{y]O�9��b5u5���W����cn�͓��A��CP�̓WMG���5a��Q4�o4r<�vu�U�	�1^��t#��g���Q�uu��4}8U�^�ʳڊ̒�f��Eؕ�@�ƍY
���֌@�]a����{� �T{m��e�]��=;��*�]����P�>��|�&�}q�����+�W.6<��.�y>���⧫��{z~��S���g�P�n�|}�����hd�g%HG���?�_���ڲ�Zv��O#�K �J9��J�*���}o$O ���s����t����ܮ��v�Gܜ���[uGIv�k��u�Һ&�}?N��3��!�q|r<Ō�W�h��稻wmo^���mٮҫn�	-6f�]ĩ��8�ٛ�^=9�gwUz��]͹v?Nw��v�߽j� ��+�+�,o42�U׃�.}�����dj:�.��5ޞ��O�Q�3��Q�?m�կ�R��i����"�^�A�׎�;Ƌ9��,4�+����e����h�wF6�읳g�Z�Z_5>b�0���Y��U�&�_���x�>BB��~�ڽZꞭ���p˭���ӓQ7��I�r�J��Fd��]@H��Rc2���������=����{G���7Dh�հ:sZ�ꞷ�/ja�ht6V�*�?�5���c�&��&+XmYcH�L*(�.zK՞�X��V���^W0ڮnW�����B��iXp"
�T�{����tǢɳ8.T�&���S��ۭ<-ϕ�B�>\�];Ҫ���S3�����k���{��/�Z/]u^Hcv�Z�^�zZZ�R�9k���ƕ1Yx�Rf��r���eMdkki�^����
�q��$��B�T/7�_����P}���Ե��蛷yh]�Z�����W#��=��V�#d�/iQ�P�v�'����9�ic�}�ߪ��[߆���`�q5�����5d�����I�6�t��Du̮��ɒ��p����-!�7V;Z�<�����>#L�J�c5��>�Œ�v^�l���{M:��� �4�Sx]}<A6�_��R����{���������7��3�ݖ�O}��p��>�{g��	���w7��S�Τ��K<i+C�Ӗ��+���(d���Î�I�	��)�E{����X�mSIAZ�q�Q.+*���L#H&<�b#C�����G��7dۚ��Zic�y����>Qp^&%�����>��>q���G����:
M/l�=k՚�G���A�:w���G�7R�N�m.X�	)d5�<y�Yg�u?�=.�f��4-W]�bڝh���64�-c�GQ1!��(FU*wH[�r�2���q��.z��n-��;oM�s�V��j:����G%"ix�]��[L��ҕg�*�V�������ݩ��M�ދ�Tk�Y�c��S�u�[L�cet� C��6�����,��"�j8�BS��j����Ӗ�@��k\ ́��9�0i�����}f��2 ��Ϡ����,>��|9�89�ugv:����V����x{�ܮ��0t!���u�7Q`iz���j�����ھ���\�-U��6��^@\\�k���Geb��^�{F��ܾ��y�t���#�bB�����C�Ok+�G�����ï~��K��-�Ϊ�\����M��e���գ�t�b�\T� u���ut��w;WL��m+Y��I�X��=(u�,�ƪY~�*�����r��y������r������O~���=����� �?���o�޳���[����̯�X���/�}K��N��g��j�����L=?X������%c�r�_�n����Q��?`@#���10t?<� �$�3nF�����.BZ�Ѥ��㖭�p2�bD�ϑI�&�(���x�FzO�+��QJIl�,�d<U��a��ve���T��7Z<� *Q�-7aC����3�0�#�V@x�����c��x����ݦ�{1�?%C���$ 䥁���S��o/3U�9�/ˍ�A2�*���|�N�ǁ,c��C��}�r�,�h�Z4��>+�
|<��:��dgǛȲ%#�&6�G!�<�>tF^Uv�#0����)���œ"cN�e3�y�d���r�#nABϾ�� ,b��	�� �M�i;qM�Ur)�,Xј�� ��v/���5�'��ȳ'��>c�~J'[V 86D�$�}1����V�"��X���ZV�sdw����
wg,d\�-�Q_kI:>=ML'���p�Ȏ�I�`U@ r`�:V�� ��S�*1�P�=dX�!Y�Xr!Q94�i�%�������]�⫓�Bk"C�9��|� �6n)R�%-�<lq���'��&KeJ�l��K��9�P��'��x#�ee�0�N�n���R��k*����
��^hw��7��qV�������%(F�%+�1M�c>aB�����l�+�Рɝ�Tgj 7ۉ	˃,gf�^�s���#'.jx#5�S�����<~@e'v2I�X�Tƃr�+dQe>!���6�Gy��g}�?Vc�G6%���+'�+����d%��Ց@&�n)̇~!�}13o��\�9��֥�M����1��6w ��c��sH�J�i`�B�;O�$`[Ш*Ӝ�*�u˝�m����%��H��u�s��)@�$��j��V1k3�\o5D�*Y��*X�_4�0nKG����-�F0-�CK�&ɩlz��F��k˃*� �tU��6߉c%M���5�Q�R�����'����:�uvݙ�Ě�ϔ�QZt�ҡ��3���8�&�Ⱥ��f����0�4����C�Q�pA��L��[� ��R�,c�����<ޭ$J������29�Fܪ��; �6�yF��jNR�C��&�U��\���J����x�Y�x8�R��^N�;�k�R<���c�c�Z%b	n;c)�F:�{X�W���f�
�}���.7GC��4
��!,c�9�"�of���uL����&���yO:n��[��~�d:_H���H����H�-��~R�� qR�0�=�݌�X�t�L:�� ��vQNb+9�#���|YXP;��á_Lda=�<fe��j�x֬hJ��U
OR|6�i�c�zU��g�-̱[lUh��Y79�'rF�/�hX�L�I7
�v��3����k,b��V��HI�6��bq�J����Y�r��/�?�`���7�Y�b��*�|w�<J4�ǽ	y<6!������YUf�X�����EVɓ��H[��%D�*�c��~�H
[e�  ��~3�2�A?�߂��dMқM���|(?$�8���1�U�-��RŌғ�7��,T3�����T�a�%�"6dq��U�Ll���\�&_
n�jG��b����`�)uvM���lr�6V����qv����EVtr�Q�R�$�VR�Q$i��l���Y�� �K��������kdWi��gr���`+�TlCS�A�O�����c$e���<��T+��d*�Do����Wp R�p��X�1 ���H�t�~;�����w;� ;�Lf!Y)�c���l�ll��Sˑ�ч��-���� �`>���Ly��у-f��m�.ӓM�Y����2Ă�������x�J����Dɡ����M�6�L��ևrʻ���Ǒw��"�#�!r�j������L,���DޱWZ>BZ��U�x�[�eX�T/9?�Y�̱��|�5,!��c�r$"�th�"�d�ׂ!r��B����d�����lz�ٔ)��|IɼS[���;�+�'�jӤ��ˤ��Ρ0���$S�V5 @濋�X�v~u�wY��Hc���P&q�%/^J	� ����9���6ؖ0��vCpFWEKO����%��f;��jw&���`�6�"֫ژ���VJ	!T�o9?�ŀ �(o�$%��2V�߄�q�̩ �auf�?q�1��ՠ��v� ;e,b����,בAU�&�̭��y�~���F@�8�cW��R���x�7�4�)��g��T1〈����@��NrxRq1Hբ���rn#GT���L��Wf�� ۻ9�`�I嗶� ���**ru����ϗ�|JJ$�#+�Lc���b�4f�4�ί��<q�#R����x�̂W�c�9�0x̥�R�K�J���Y�y��)y rT�pV��OĖMQ��x�˽*�+�I�Vh!�p�7���&T`G�� �]�s�#�%2�$5i��,8Ȳ��]�x��U����)�ӬD˧9���WڹR���� u�2����d2�V�L���a���l�	'���$M���2@^C0A�Ğ��+$fug��6a�:�"%?��ƍ��B�d��T��;h.#���J�M1�T]�$	�*Q�ٸ)��,}���d���K�=�Ra{|���tŕ:��5���:C��!�1�@�S�޷��}A1-:;Ϝ�e{G
l�d-fP���uZ��m[�K4/6�~�3i�w�Y�g����V��`S0=KyIj��c��v�Z-�REJ4%`
�����e����G�`V�����S���W�N�띎���8�E�z^���ms��yԚ�'�||~����;Q���*���+���Yz��θ�4�v���mޘ���7x�C�]���)�e6(C+�[\�V9����"J��Sk�li�u}���(#�"}N�<�\r�T�1-�5ds�&�!U߱\��ws:#����۾��5]?��)՝I�:�F�M��72
?�a�e�Z�V".=qy�R��1Oȕ�>.к�jk/����F�F�H�S��<�)�9W��$Dx��ux�8�zrU�=ۢ%��I��¸�.�E�&h�WJI2�=��:7ڿ�w�=u։ԝ������Lӵ�7���F���M4�mP�}��\C7�O�tf���iz�c����ֱt��2K<���>�Яs�[��M�4�?g鐝B���b��9�G�|SG�=h,��֖N�F�͸:�z]fm��MX�k��Q��x�-Ț��p�}���i�Dd-�N�����]��\wGC�Wb�á�����*���O]�9ʘ8������Ȟ���Ԥz���_Zbe���I(]����S4-��n�n�l]Q�c;s^�:2M<f)R}QY:�ݫ��]s�����\V�}A�:���:����+�[�Y�W�Y�ܣw�M���1y�I=X��uh�+#���q� M��}���QGJ�I��n��-+���=#�n�wKE�4,M���������������l���Qbj��	�u��d��o�;�n��h3؃Zk�uzr��Pe���nPö]�D�*�G6v��&�SE��������U��"��2pY
<��k]��i�f$V�僃�z�M�r鮥���N��ޭ�n�bǡ���s���_�on�P5GZdt��zm��w�ky><_��	`���F]�?��ZO�v�*�lj'��:��Z?���܌E��<��}�`
��N�a�#�Ԭ#�VԺ�[si�+Y��(�Q�=�T��� 2ݩ��V�<���
�ӽ�^sB��۟}����W���K�� ���w�����Z�:�D�e���bt�]�6����#��t|Hi�� ���z�9���C�Uے�/X�-�v~�T�V��ۅm�"�fqV!�,�%�1�̪�a�c�oQ:�퇩�Դ�G[�Z~хf��w�U�S�,��yJ�<$��,\I��g��p���t�����h>��{���nWq����_��+G�gQ��������K6���gU��ɑ�xz50���m���e��VkM�`�gJw�����>ԜE�$f=�`	?`� �I�"w�C�F��	��'�.v�Z8�JC�D��8Uhde#0�;�Խ����tV���{����_�&6Fd=�v���'��]W�`t�u1���
��g9zv���|K� ��<TH�ǭ>�ӓ�[R��;������H�۞t/YL�2ՍC�XY����c�����M�5>��,�iԥ�%`�~��{6ƃ�h�WIe�`:Eqƹ��ۖ��G����]�=C���t��X��{zL՟N����kOMÑ���4���3+���'\K��8��_zwX#�c�#mP��n�6��q�R�G���ykXyX���"M��yS����u��R�t�w>���i;�Cޠl�V�[RSGiaYb�ȅ�e�'GY<R G-��՟�/����<�����ۧU��3\���w�o�]Y��=I��8~��{o�����[�Tif�-M��Z3կ_� -��ܓ�f�F����`�����J���gt������#=I����-hQۖ�Q��[^$�E�;��j4@xH��1�
�� {�t�k{�ؕ�TT��-{���\�l�!����'J��~���~���N�?�F�i��k��q�lF�����Ȇ/�k�_��Qt��q�і7�vxE���ب�[�x�
h���Q�C
Y���tWV�øz��i5Q�i����(СJ�W���jG�㺅V�O�I{
�o�f=�����������׵�t�4%�t����]8��q�l�`���;+�/JΓ����/�'�#�O�~������ּ;�f��iڍi��Z�QjRX%�D6� ��G(C��W~
��Mj.���m��t���z���lш��ن��EI�ˣ�U���x�tg�c����3��i�u����>����uwe`5=3J��u~~VN����,};�<?}N�D�ԟ��>�j�7n��bׯ����l�n�W��4Q�����d�����_⃨Zrm=�F�Tx��d^��t���m!�C���]qoqF��מ�����>�Ի�f���潓�Q�N��Jh�n/Ch����8&	ѽ�����M2}a|ZTg�Ҵb����>��r����=��*O ��|��5�G��j���'�4�		��D�zUMP뺕�����:�؊12�
��T�G!n`�������Ϟ?H�/i�����ԗ����A�Ȗ����ǪqsF;Ժ+��2�]����]7:2դ�(�fx�֗K[���4�n�����ڪ�$��+������F9�:� ����.`��z�E>H�O�RP��,}��͕��_��gZ��M{��������BǨ�.����4��_p�a��f�Zu5D�ȶ���^�O���AƗ�e�T��ؘIh���Ix�,H�W����Q�G�d�!s��2�Q��T
�G�)������!�8C���������W^k���t�.B�������3�Η�Y��c��q��:��4#�h���� ��ez���e<rY���nO<��g��灟rMX�;{@���9$�ϡ��߃�����~�}�i����sT������g�u�u�\���~��p釋�h�?�F�jt�[P��&8�1�^`������z$숬s������f �pc��#	+���<e��U��I���<��j�o�8�ȑ{���#^���]�C��M��WP�S��?V�:���W�R�pM�t�,�CM�)�=������%R �Z+���	*y��GU�!pce��!��C0�)>���SK�d�lx۴_캏��9��H v����3z�!����t��Gw���-���ӹ�������8��1��nTvz�n	�]6��:�F�:�
�{��/B@>]?�	��2(#��=���}��Qip�#I7�`����	�8���s�^�����>_Y��5.���F!s��j���I�ڑ�I���������i�"la�[�%O����� �� L�v�؏�}���?ǟg<5o����0Um�Է&�نa�}� �=V-D��@�����������i�v	�p?o�����l��g`��%��o�`�� ���z�z�(�ny)� ���������q w���Ƴ8^M�7�lXC5����Y��`�D���a��^uu RO�`���@S�oh���������}HЯr��?�}� ��� �z^�ҳ�fwƠJf	�O�V��)UX�(��c��~�����p��z��r�� �<���X�<�|������� 1��C�O�-�mB��8���|<wU,22(�H����n=xOZ
IeQ��hn���� /y����	*���� ��>���k΋��������Ǖ$ٕʨ����X�P��^-��bJ��PG�v=sY���G{/���?�~=�����pT+#�>��?�p8���Mk�]�:�Lj:���_�%�j=��:{5���|N�ճ1����]R�c-���IԤ����uF��Z:�i�/c�]{x�cp���s� ��o�ķ%��0=�:O��V���S Pξb�"��W^�;������׸^����o��o���}�����M��e�tΫ�9��]:y��9�;����g�?Z�S����O	�c��tn��k�m�ٝ�ƕ�k������5��"�Kd]�
�4���V!Ҵ�̏��;�ƺ�P5�SI�om\2MV�P~Ӣ���:9��=�a/]Ӄ��觼1�r{u�Aw������s;��[�4.���.�df���Om:wJ��-E:G/�,���gO)%9�~y��¢�p|Pu7Nܚ���;���Ѷ��Ub��R�"Gnx��l܏��ox!�+�TfoG6dt7n�}��n�����ӭ+�Z���Y%��I9�H#�k��H�U��w}���g����w��K�,.��ײ�eԷ�Or�5�u^F���d�\5W'	��D���bz�J��)L7�XH=#�p|C�ۻdu=t��_O�Tm��`�BCM�W�ri�t�n��é�jס��K4�ݹu7kX�Z^�ә%��ۊ�h�fy��J߼Ѭ�{�|��"Z��՝s��^㒻��K�O���
��~�]yԝ?�j�;�'�]��azӤ����^�{�ګfe
`O%���hy�Z�����dn&.��2l��k���*���R��Xܲ��5:Ӥr�m�;Q(K�r�ee�� �/��Z��*��}^�.^�䭠��U�xuB�(Y�BRY���{�%���d��:�U�ٷD���������n�uEj�a��##ڎ�v��t��.��M�g�Z9�˞NiԞ���u#���a��{iiM{i���bx�'��X��ޏ�=�j#��$�c*-x9�Εt�cu7fi{�^�SYY!�E�:�lx{��(�*����8S��O曼q��tD�.���=����{��^��ѱ�S��ڿlu�_D�[=u=C�q�<�Y���^+�i�p�ǫo�oR��V�k{{$��g�|�dMY��/]�XI'��ñH��&���+s�� ])�}3�.��V��[�B�V8ni|YV֖*�`�h�_#��*��s+��9����}�wӢ��-/�Ou;���!���/��zG��,}oH�-;uƋ<e��/Kȼ�=� ?X����=!����"�>��t�R���Yw��_(?C�l� �/$Y�R��2HG#H�W�Ӹ4������j���<D��x�`T�Z��<p߼���U;��9�Y�K�]�����o����>������tA��k�A���q1��XX9�1�(�7�|�#%���LɄ��W�k�1u3[�5}��)S��z�f�NT��EY"X
?�%Ŕ��A9����tN�h�h����"@���܅��Mfkl�,����7��G����WZ�Q�:����7����k��u~��.����+�:�Z���ԡ���bt�`�6`ѓN̠7�t쌴�9�Ld�ρ���m٪��w5	�l�zu�u:7CY�NUh�P��2,-`�X�9fO��M����9��+��J�E�4�B�zN�[��l܌K�-�k��Y�?v�:�x~<u�r����H�}���s�A�z,�՚�tr:b�S�ɦ���u�.�k�9qm���~��tgJՁۚvܥ���~U4�eX���������9����oԴY�[��5���� 7&���{y�����O g>�:׭;�{p�?I�������J�q�MW��:�M��r������P3!�?/'Q\��dC��������u2�z��r���o5�vd.�%�1$��4Ů 0|�(�΅є.ws�P�<k=7���^���C�$O�O:��b�����E�o�9�tw1���kZ�U�2��ޕ�-?��:��'Mv��N��x=*�y':�M>��.�IlE�$i����F§%��_��:�5;:���g>�j��c�<÷��<����<������(�� H�D�M}lX��{��MMP�n����R?JBfU2�b�FYX��'H��,�<>�u�RW&���tw[R��P\�l��ҵ��2�S������Oɧ�A���T����)�v����EB�����>�h�:��S��~j��{Y���_:?�����ɨ]��0C_FkR�n��Qs���!x������|��M�_u�Խ_�z�{t�v~�����_Q�.�Ա1���A�J���c�d[;S��q1ޘ�?��D7>on6���S[�5�sR����c#�#8g>S��`��� �@ΉSЫ��h�h(��\B8j�E�:� "B�U�W�H�v,I�]�?x���}yܟq�����_X�k����j-����5���D�1��V]�꼫տG�ֶqT��_^ͩ�h�+�}h�,R�	S��P�������ퟫN�Ҷ[�������7����k"�'�}���K�Y�����'����^����ӽG܃�c����G"���^���l����PƎ24�d���O�;0�~'�H�yZh�Au��2 	=���O�_� ˔a�������I�1_�og���f�{D�>����9=���3{a��q�u�g�Z���\L�31��������>���D��E��jm��l=���>���s�����G<}�-��r@?�@~A�����_����~��t�v����j]��7�z���ǐa�]Y��F��i�Yu���⾄��Q��q���gW)˨i4�8摥��	��cB�������UR\�I>�e���}+�gN�1�(���W� s�a/s�=�=_V�z?%z��g·Q��9�/:�ɞB���,�����l�;Mp�
�<�+"Q��J��4�)U�B�k!$s�I?��I�{GՕkذ�D��C�>� ��J����r����Ӟ۶~�{Q��׻wѝY�uw[t_Ka��w��|�N���g�'Iаz�dxz���B��OW�0���L쪥�񖅑����`�Ͽ��y�\{˸ub <�9�_~3:B�������)q�NYfʊ�J*5G%c*m�Q	���Ϭm|׫-9�)�.@�Ӊ�d�`Er@w}�}1c���(f���+?��@l; '�&@��Ţ�*�Z.q�K�N9��Y��KD��U���D�|������@�9E ��,���M�A�0��6���pC�6B�ZV��tLyŃViWV�dO�14��V黯%*~	,�������~)E�^A���R��d�_8+��l�m��Jc*Q-�@���ni)0T���BΥYv%�p��-��V\
-�����I.�5�P�%7,y��[�J�δ��x�7,̙�S��wDM����r���I��R�Im��"b�s���K�R�_e�E`�UK��ے�vBVE�3i)(�5�2���P�v�j��0a�T��j�2_�v�O�Tl�j�D�j�_�Q�f�9Y�,X�(+�NT�8J�^E��d�Z�j����J@wO�M;�+iTR�D���d��M���RIG@
�mTWc#0�26Q;��N2gjV^P]O⇒U��%���B@����%��Wa�9���̙�L��N�>G졷$�O2]dJ�)c���v�(��QH��{�ʌ�C�%Pf*�`]��&�4l�R��Wtk!O&<
��|R�A��1VN�2 _ Ȏm�YL� !9'b��Uh����v�e1����TDeV�+cNu,����ŉISy"����>���Ѫ�ճrNI`����n�V-�u�~��6�7 �23_|m+1���Ґ�43�$��U�|��]�,Ś�ES>1Vj�责o)HTY���9%�ԫ~�#�� ��*Mc���|�9-Wű�P��1��x��|(X3`BzcļԾ?	�����Qj��r4��9�� ���۫I��Pϰ�A�f"�����(_.>�B����X��0YYc�0�RZ� �S���9��_�8��M�_`J�|��Eh����X�O:��O�_��$j��#"˳n%���D��R�l������d�<b�����o>D3���EѤ�5E�'EM"�F6Ev�曞G�ݕ��c)<<,cX�c��Ňӕ���J��$�%@vfVf1R�U����UAt_,��i�TRSy���*�� �zc&ϒ&�G�U�y���t�,���X/��ᚊ $,c|�<�^Y,�x���$�\`DY��)5�O5S3�a*a��+7��LnHD�����b���5��~��R	%�##�%i���e*T��ez�
/n@((T�Ա�\"eW�PJ90�(�{�G�,�WuW��<G-���k�'�4k!��!Y�m�N�/�+O�컳6���`������v�͚b�����WB@��?R�N_bU�1��|e�!��P����J�p�s3!��d���1�,���3J�6jU�(�ڮ2*���bH����<}1�iM������x9آ-��,A� �Ua�ĳwF1�$�NR��[�+�ffo/ 
)��ٛtA�\+1�q��jVyUf1��,�bb�S#�f����;�r}1��dA���b�yXddη�ٝJ$��Vp��  o��Ǒ��R�Hʳ�j��eR)�*�IΑjP�5
	�������[��\�g�fbY��8��H�H��I� �}1�ˊT��	}�$��C�c���7�Q��R��
�óX^����͞j�*����Jd�bDK}2�(�,eXG��٫I����~�<rQ~B��@Z��/�Ee ��`M�p�.;��� *�Z!�+��  ��a��L������d�Y�Xt�9#�rQS�-M��37�"B|�m��`%,XY!H�C�%.C�!9��$W�G��}�7<Iu,e�Ch�2���&Մ��T�Dw�DP��m����d����U(&���f�(�x�J��%���$vm���HO�0��H��3[�ڦMr�0H��G3)؏�U-9��A>���?�qi�4�XL��6^&�rj<`�5C�@�L�rX���2s���0Z= ��m��{�υ�M�k��Brd��\z����<G�'�/2�%B�&�*�B�į�nY���%�>E�q��j�yd�&���!c��T(�c�t�G
Y&�Pp"O��/1��9r]�r� ��s*X�|j�d9)�P�$f�36"�ɖ\ (��Ց�^D���$��ɖ-�j��3����?##�_�q�RK�c��k�ո7�awY�nYQ�M�a���d ��$ٌI�>�W�V���^O��ъ���Y_�7.2p��c���xK~G4�x�^�$��?�гr'�h̫�n��������tZOuiʲ`�	�(,�9���f���P�22WW�B����edv��o�,�d�� Pw(W������<���1���?��>�3TڛqFf'rG2v.3O#M��5�G'E��qq�;?U�uo6�����uZ�y$�a,�Y�(]���t]V�7�Mѩ5�eF
UR(c�؞W+z�(--��!�G.�-zƵ��[Q�/%
a�%g�&���1�2ObV�b�yec�!��연r��WE�����~��O�+�������-���?Yt΋�\�J��At���Z��e���ioE�ҭ����o����FXlW�џR۰�-�p�].��݊�׋��"��L#J�S�=冾�]+���Z�~cSj:��A�O���G�rV�������#�7W7��OtG��{c�� u�h0;-���[j]���|:��p�~�M{2�g�[���CY��kX��Ҳ�E�����|Kh�믛�Eݚ>�_C�5DZ���CԌUE[��6"�U�q5+RH��GY/��M�ЊZƂ�d��뽫M�#���n�ݎS��� 1���f�ګ�dl懴��{_�.��a��P~��WTuk�Z�έ�:;^�C���-�Y�mНe�R����kZ�l�f<��;5 �鍏[^��]�G5M�ԝ����tM��~��igC=h�v{�t�>p����DF�'Թ.����VX��gW�꺭	(ƒ����d��q��z��A^�$���)nu_�>�z�ڧx���ܽ����[�=;�]~���uӝҹ��^��V�ާN��GY���)�=6��%ؖ4�h�����K��x�J��N������{Z���AwO,���4���4$@�O-!#�xGp��������~M2�ocJ|kCZ�a�Yge6�A/��q��x.��ǒH��D�}i샵�}�n��˧z｝�ǞF's:��y8��K��BƇR�P>O[��5�7���]~YOn��[3*��ZƏ��1K�־�j�f�tN��ӣ����)�MN?<;^ܺ}w�2I�m�	t�B���~j�|mْ_Gz�S�2�#U۷�rA5�� ��5yu�K��m:��:��F�L�[�8�!��G�j�ϻC��k��Q�Ow{y����n��Π�Eh�n�o��i�����(dg>���K]���i��]K>��> �kF���ҭ�Wun�{KևM�� ҭOkO�$ �kZ�D�������-���$��G�:�H���*i�3�{􊯨A6�L#�;N�$����ax��$-nM߾�5�};�#��~�{���#'#W�.PuX�����\j��~���m[_��y�S'�1�iS��\�H�t_���s}չ6}����@T�r�RbV/Je�c1���1���d.X����j����i����"�N���hV��Ւu!�׀�8FxԮ�mُC��7�	�N��h;L�G`;��ϭ0�O�#����.��W����մ����P�f�d�W>�a��h2ɽD�v�QT�gL�t�'vE٧����Ff�YaD�;43
��d�K��r(�Ubb���}��������J��v�%�Rx�)����쟼���]��5yÑ$�:�{_n�����=w�w�{�� ���^�2:/�������~�N�ˎnWQCD�:{OM/��Yi�Z��Z<��hc>W�����c�&�U����K���CO�c�Ŋ΂�K$�d����b�I
�e�.�~|a�4�F��N�73IN+'���7�ʑ��Z�$�9��q�4p�	Ǫ�����ݖ���K���{����=S;���]��j����N��i,-kG���C�b�jq�Hɡ���d�?��?��YԵ�4tG�S�7��/�E��"*�]�N���Q+,r�;�=�O�W�uK����@�^JUL���*�,��$�#�Q�k�f����雦���-��������b]���uf�������2S//Bִt˦����]�)�� =뉕8��ⴁ��o��:W��U�cc�mL(�0�X�ʰ/�X�$�!��1*:3F�QK㍄9[�]B�'�D���s�����,�V�>�ܯ*�X���Vc�$M#-�Z	T�;��ܦg��[��_n���E���u�V=��]Z����N��ҵO�k�Ԛ�B��hPԒ8���llF�ޫ�/���|3m��F����ͳ�k�h�1�ue�Fü�f��f��� �x�:HG�W���?�>���:��k;���ZO<��I^in|�Q�V�=x���m#Y��u�B��޻��{p����^��~���N����H�β�1I��.��r������-3)Cx��rG��� �3���j�R-"�3��zROA�L/�f{3�^6�B�$�R	�=�:��ښ~�cM:�۵�ϪX���2��^�t�2#	V&�!{�����Ӹ_����o�A�~�������N�����N���������l|_Ǯ6S����+3��$3gj��i;+���GU�����ѷ>Ж:�/�hҴ�h,���"x�g��XҶ<.�5#rn�� ��+N�n�.���W��z��VȔW�yj=y�f>"��D���<��6��g��U�� �Vt�f���︰�~��_m}��ֺ�O�yڽ��
d��z-�_u�L�R[ʌq9�
C�t�:���!Lkz��^Q�����{�L�Q-���1Y��H���ȳ�:�W���G�w����h�~ȢgmB�2� �j7$�4��HYk�1�"1K����� Lb�z;���]�����u�Ih�E۾���2�1��OP�����,*�WS��Ķ}u� ��8ט�~O�\��^����nݷ�Mos<��Ն1��9>m�d��xx|.xE��\���4����*�u�!X|24l�]T�2K��T' �2s�F}�{,Ӻ/B=��;�����sR�ѭ��gq�������zc�~A� ��Dr;��Z��+����7mF+�q����7>���(\���G=���ʕa Nc�1��Q�{}���k���Bm�ge�<�Gp � � �_��G���_��1q��c����uN�Ճ'����Y�==_���OmC�)�y2;��h�l-1ej�_R�f��Sڻ5��g<��F>ô(R�I�-�"�}Ǽ0��P��b}(<��x�U��������J~�v[;F���ckZ���պWڷJg�7Q�ְ��Xa�?_�Ξ#O�vU�D��Qf�Y��
�=m=k(�H~Þ[��A=�p��O� x�$���,L����C�-�A�T�x�<��{#��辏�yڎ���Ww��������L�z/lz^��e��:�F�����E*%�&��#���8�tr~]���o�>������ *��xA-����E�p{�{�"�P�y � �#��a�=����N���ݶN��n���b�]��MG^��L��)����f��;>Ox:�V|\KN1T��3���Y��-YQ�Z#�B6N�Ok4��U�ل�����O�=-i+7��W��9`œ�Ujcb��P�Þ=rm=�����v�{	�9��@�GO��E�=k��w����#���N�y���=3j�!΅�1Ǭ�k�[4�^�����'��n����>����n9��H�\��F�@�5�'�. '���}�����	%)Nqa"���� h�w� ��  ��$��$��oǳ�������TT(,����lg~r�D����C�����$�^w.O�n}U�������}��9��J�!G r}��|��墼�'*��ī$�
(��\�l�Q��~w�?��Kj͊_��S��~G����9�C`���z���`b��\O����o�� �L�����_0�SH����'�}� ?����J��:���z�}����s(a�6��izve�4�ye'����0��C�́�~��v��sh�Gb$
�}�*����}���:���1^W������?'���������6=4|���ڸ�������L���(A�D �W}��X�]BΟ$T���1��?�x��������O���-��xP�s�������ǣd�cL�u��,-24�Ȧ�6����j��T��,�}�/տɣM˨$����Z�p�`S�G��?s��8?|��F�2<��J���7$�$��G�l׵����5�K��c�?D�����x��I��_�����)�=;�w�دKu����q��9i63eMA*�)>���.-�>�6�����V�ȿ2"�X�
��*����G�<E��Q�H��u��#Ԃ��=x�V#��\+D{xHhC}2������ �N���� p�}��R�l2k�z/r3:�[��� �h�����g�K�05[�T���[��D�5���=!�Ƭ1�}����~�t�G�gJ&�{W}Mt� '�Nգ��K1mr��9j��"֠ƲK4��8^[�i���&�SsJ��i�IhFb����X�2ҁ3<�g���s	S�[��#��c/ݗLv��w��p��z�Q��L�t�~�e���v�M[��ܞ�66f&gOR�h�4�R��G�|]A�e�9>):�~)F���n��/6�H�L�"�#�^cܢkM提�)<=j� [�3)4�WO�Y�R��\!���3D��&@ѬR��h]9\뾀5��a{���QW�>���j=U���躃����d}[�텓����ۯ-?�4�H����J�|��7�eb�>E�4��C�%��oM��sa� \5N�ֆc���z�U�<fXu*_U�7�"b�V��k��l:�d���@���w�ʏv�"�Ζ@75�>A�r�[�|�·�&����º�T�L��i>�:�w~���]��z� �4��vs������=7A�^����qq5n���ѝ#����w��DZ��	�&���MGPĜ-OU�l閡����:NЫ�˨ߊ�zr=�zTB)�E>�5��Mb��֮m���ؤrD�>�u6�Ww��grIv�U���kM~u�^(+�i���Z�����T�q#f�{g��~��􇶞���y��}���.�״�'��;��=>��W�:ϸ=}��8��֣9�����,�șC����	�Hٿ]X�W�]���vk��0�Zz�"�hIʽp�Fc�I
����;�ᯥU6��:���ڍ�ϛO���5#sdM"��T�G>��j�{=�w����-ߏk�ս��7�;KНw��t���Ѵܜ�LmGQ�o���vT1�L��d��ǭi�i�
ߛ���-����ӝ��.���N��uzj�&�/�Y!I�����#D�3�N��8�<�q����ʹ�c�-�أ2�t�u�V�C�CJ���IZ/s���W���0R��=�j]Yup=_�vǨ��ۇKww�N@w#�N~/����r� ��|�\`lt����|��'�}`�^�G�%�~ߋGu�� �.��?-3�W�9�$�eR�]g>0�<��s ��K��W�$�֯6�C7��ԑ��Gb�ΑR�V�*�4����ӿ�x��k�R������{��8:w�{J�X�u�j=���Ί��!̬u.���>���q�Lf�}AqE�N)��rduG�������=Id`dx�P�f��t�O'��GI;���}�g`7���%-�?�=Z+�ǁj֖��@��$A�,����">��g7�������w����V�|�N���ˮ���ص��϶��XɮC�:����F�sqSV���^�SP��Ro�݃�����en^�h�E�fZ�I�u�%�j�,'�O�z�9�~%���J�W�s�к��6�L5V�����t	쯊Ɂ>ef������/+��P��foC�L}3O�����S�;]n��O���}��/�:�P�]�܏���3#;�X����m<��ӵ<l<��θQl��jb5}�O�(|���=;N�D�\V��\���j?5����A��o�dQ|�-d���KU��WM���V6R�(�Q	�k��#>P��	n��߬� V��D�}�?��jYZN[�oS���g��B��|�ͯJ�Xxyǧ��q�̹�o]Bf��8���~�j;�*օ4U�uR>F(�%�ح!��X��L��P�g$���
���-��5emJ(ݢ5��ԑ�������i����# ���tzv��^�;٪{1����SS�i�>�љگNt��i��i�ڦ�Yc����Kb�X���x�6��]�����э�k�W�]�Z�1�u#����AV1Y��-�_ĳ�Օ��v��:�P�߼�t��@���I�����rCj.�"������ ��x��������~�u����=��WQa�GP�}S�q�M'E�.D�~���H���.����=�\��A��M־��Gv��4�v�¨டalNS�I{�(�'���$ eq�7��[o��k����>� ��S���� O~���f^,H��0��3�����).��7v����wc�:��]K�Ԛε]7�zs��?�6�:nNl�+f�����f3C��_�:bM�Jڦ���옡�/��E�B�L�+q�)<� ���z�;�KTV��������#)��n8<�^����}�uǴ������K�z���l|���GRLZw���\�gy�yM�zo��yH��yCq&DƬ�'m�&�3KD���xO㰂�s�o`�鲮�y�Fs�ϣ�+s�?R� 5$�8㏱�7w}�w�݇U��H&�i�څt~�v;�=.�?A�]u��WI��@�p!�\�I���j��9%*�(�#P8�8�����������K��O�{'�7��������ѝ��oҋ�n�k�l����<w�;e (@׿�٘���_�_[a�~��it���L����媒�N��ʰK ��Y�bC2��@?��{?���+He�w�*�� �ow���9�r9Ϊ����i{t�uܾ�׻�ՙ�e�{O��C�t���lXh:�o�#�4;P�].��Q��J����9էXby�>�!z�c�B���@8��/�иp{J���<�=ILv]�34c�7x�a�/�(A���x �6����û��&��ks�k��N�gJ�8zRgu5%����j��i�)�̈i���fi����=%��Qn�LO�e?o�ё��H��c� ;��t�
��
����py�#p{��y �8�8Yܯr�џ��n��h;�c�?���=�����]w��u�)�y(Eg�`}�Q��\~���y0;C3��G�s����¯.}��������?�t�\ɡ�}$ʹ���1�AvH��u��-M�ӊ��o0��3� �� �� �����?���s�j>YVw[�,�Ǳ���'GC#F�!|��`�K �v��|�7����M���#LrV��?)�2ɐ=U�Ve�`X�|��Lb�I*V�|��h���y���Sİ䍘�x��l�Sc8��Z�*����-��O/+���Ā+�c#�*�y"�Ik�t��п�dN�\�q�2��nD�Pb�v��3�Zm1�����3٦%�+=�䱍�dO�#�B�"���x�6:oU!	���v���˚�����h�gjboO��.7��5Bq(ޘ�8z�I�pg�XeZI�uj�o�xY�F���@>=1���'��m�u���u���~-y�8�Ȍ\�����|=1�2��HT?�񱧔�[�+d�mL��ꡢ�ɿ&��geŬ؟Zaʘ�>~)��D�єp;��!U�,`&��v���g7��*o��ơ���c@�<l��Y(dʜ�����NBF��b�֪�j jD��Sf1�mL���I���6zL���Qb#)+ʖߚ�',�'�B�>�GǺc,+��e����9뻷 �U���O+�LKOl�b�ec*�q�,�Q�?,`�
�V5\�^	��.t��e"��,H,�ID��(QF0��T[c,d<M��S.V����Ũ��ln�9�R�C�Y�j2~VDI���y\Q��ۇ�i���1�Tc���O]�0�5��a�ǅ�����Ǳc	��IÌ��zR_d��)d=�q��u�PX�^���g��ql��hG	c�ڶ�SY=m/�����`�1�kJb���D�;$��ř�#�y�*��C?/�^{��5��8�g��]���ʅ�	Gr) ]Dуә0Z�N�e!�ֆ�=�������y���EeR�UO�x'�0��.ge]�2	N0��$�9�H�U�SdC�ynAo�c+����#3:V~*�F�~,��E�����e'�JD��z��3	FܨV�9�,<Sȣ*��Aد�1��<�6=�m<�YqJR��8�n"��<[�Y�c*X��l3�3������6V��v��x�ӈ�Lc�&���Ş����F�<I����R��Tl�R�0�OǭJH�&��]q�$���1k��z �P�!��:p*�+>h�*#W[�q2)>E�ꀉ�b����u��H��?"��2�r�>R�3hc���n>��@�0k��Lc8-UQ�JZ�B��;Q�A7+hJi!,9 �X��x��T�)j�d�h��J�7� �!���Dn\XǼ��Y��fɬ��o,�0�f��"1b�Q�\1��l{�P�W��V+J�r�E��V��pY�NHX�0�E��Jst�����ǘ�0\�ra�Q��<��c�#����/���*��3�b��#��ʀ��[�"���6�ʗ~Ԋ�DX\�-X��n���i/��rܳU�G��L�p�71k-^��7YҊ��y�!	FA���PX��$i�fS�s�,�HR�{xs���nA��)n~P�ጘ1����W�@�1C� ��~Dݕ7)Euq�n뿦2%����֖um�<n�
U�����������epClq)ϑ+6�˛�U��)
���X���O�0��Si���՜2��:���	�� >��W�X@~#
�9iR&�T�K�/^(C)p�Ӊ]�ؖ1�5Z6-iIͱ��#)�+ +~�J9d$�QK���V��ɯ��^�',��DeIC�F�X�Ne.� T��1���|bt.�刾=x�/ާL�/o�>@�����Ǣҭ��w�D�[c�&��IP�(Ŧ-�	qȷ�2�:�dE��� ���L��5�N%���*�<�%��1�����&��ldzp�i&ǽB��d�%B��p�������rC~+VY�C-a��!h��'?��%���'/��tl���v��F*�~�Қ������()����
�c���;Kf�klP���β�4v�ý[�r��̼wa���h� Yyh�T��tc`�H���M��+,��3rc�g�ў�h�Ͳ(����Y��;ߑ!��Ă����Ő�$J"�bQ�fׯ��^�2�}I��1�R��4恉w��	�y($��$��� Ӑ�Ac��qW�)�3dEmm��Zr�K>���I~I ��=�i,{+-B�t�];�>��ɰ�.,�� n���jY�5q�<�K�w�j�p<�8ʮh̹�*]@*��X�2r˳��b�,��ș�ܱt�,�B�P_`�%�e�^$��E���SĠ��e������	�~)�|���1�-�.o�rS�)�c>F8gwdo�RH �پX£ֹ�Ea��<�>6_��>72��m���f^�`���\mA{��W�v��Z������z�dCO_�W(@f��{��##4M��y9��t������_��mˁe��y�jw��K��r)v��(�mj�����{��5�+a���m�Q�R�v"�N�7�V��n�2���e�a:����F������?sz7P�ot�u��A�t�g��ws{�:�Q�-�Ӫ�C��N���Ze�U��:u!4�޴2��եTڛϦ�9���[��2�t��4Z�-��n�M�>��gT�#�;�1�m-KSܛC��N��wsl�[�x�۲�����!��4�Ӊ"��E�R9e�{$]T�w��t��8u��/�s��i���έܝ�5��u"��H�s���S��/���j�)�c�$��<�&��Ü+�in��D���t�&��Z�鲲�e	o���B]g�Q0W��P����s7��Jzw�nn=2�{Q��3Sxk���+VS(oR2���V,��A��w����[�g�^���������v�B�����o�޳�����K�m�鏋��C��?4M�31��@�L�xϧt�)�l鮩������û,�R�Uc�*��a�SIZ*������3� h�;swV^��E��t�lM�t-����y�X%�a�y���'�xAt���"eO���;B�i�{l��ꮋ����3ۮ��n�ζN��g�PS\�p�3t��R�yz+��� V�3�)�Z`̖%��g���C��t���׺EӝT��w�*����ڊH���cBԫ�47�J�;�f����a.L�lMWjkz7Qz��Џul��rmsH��p�f��\��&
#��MB�H�ȫ1�xc��9~���=�v������s��h}3�^���VH��K�,.����蝼�	���ml��R�&�8�Ǒ2�Q57�_}J޺���-ՠ\:sγé\�SS�b��4��m�"�y�-��I�f�nύ]�����5���+@�ni��cL��X���VVuQ+D����*�f�{����=)ڟs������>���-�_�X��f�@vf��:�Y�����ڦ�\E�^>T�V���f�S���n���MO���lǸ(�=�GM��-سqURw�i�O���?��*�b�}�P}]��[�`A�O=�)�]���N�$�8��K4mq-�n	',�D�-i;c�3���v���Yݮ����?^vI����nP�g_�]���>��{��v�\>�tHӆ�����C�\l|k�i���Jy(��l�S׺_�t�[G�xP��������3X���]Qe�'��%��)�P�z�M��ӆ�wv�����u ��V����U�Y�5;?�����E��I�FI!�i��G��v�'nu�/s=�ܿ|{m܎����#�;7����}���UuM�u�l��i�?�>�\�V�M��j������e�2���|��뵡��A���L�}Yӧ�Y�1'����(OrMVԀ�^�A�ġ��8u]gW�(���Z���X�j��F"X�)�O���+uQ����2�����_�#Cѽ�{��� N�>�Ï���/��o�3E������;7+@�,|���������
ңN��	��֎�|�Qt�nDۯw_�n꺆�#A[�:/��I+��,n ��Uk�y촒�}�ӽ�񍨶���t䖵
�dsi��+�3�w[w���KOaL0�X�B}7i��vo�p:�ݿ�m�]�v=�Z�a�]��@��v�p�u�ό��vjn��i}A$_�3f����*}}��}����]@ڕ,��,:\�4���-K!_�+Y"v��I�\��,�$Up>w����+Ż6��oO��ifԪG~:�Cej��4q�b�<%�h���D�7hÇ�#����C�}gn�u��c�s���P��z�����t��N�^����鍋l���ɍ�ˑQ��{�
��O���T��Դ��r����^�ȱ�Hdn��pr\vđ?L(��Y���n�A��Юm��Ii�;Kv$aVF�-�P�����0J@���>�폹.ˏ�7�N�WRi=��MN]��e;%i3]#X�4�+E��ϣ�*_S�uې��os33Ӕ����޽h?ӥ�;��mJY�{��D-߿�MUl �SDw�Ȃ�6nY�&�ַ�f�o{>->���՗�iңV�C,�'a5�in3��Y_���vƗ��{Y�a�އ�qߦ�_w�����˥ew#D�Zj)�}�'@MT�OL���S�Ƴ����d��!S7M�G&�zW�u.��[�0�M_N�j�Eiێ+�c��s��O�
p���I�y�z��O�t����ԥ�۳KY/i���{Q|�H����/����I���|sG�L��;�"�~�k��~��C�g\�oL<�w�\��*_��,^8�O�
꿏�k�H��g�Qe8�w�\멿� }.��ݺΫ~�����_K�kKr܀�|Ha���nY��}��I��zS�I�C�M%6��R��]$Xl_�\��T#���Z�9sV�^�IX2H�]�����m��~��}U�+���5]C3[���OFN���v&�N�`�
˥p��SN���X��Ԯ�[Q��M���I��:gn���H��̥)��KbQ
���Hjv�Y8c��}��ۢm��5��)�;�Fa��BW�8�yMjcb�uB|�� �%���K9f�u?j�;�3�u���u�v�z�ڧS�� W�ugJ��s/����Q�{�����.�ZmZh���,�F �{n��u]1�,r�/�ŉ
�	j��ɂۂђ9'?�J��Q�A)�$d^>�8�� q�! ?P_C9�ήҽ�uS/�^����t�G�OH{l�������$<��2���7Ǎ:m�5��z|�d�Kŗ�i�D4��w���l3Z��}�����hu%������8�#��M:���k�VP�ı%})�$���s�c^���޿��Y�m+�����Q�m[F�H�/��ִ=C+�4m3���U��8���z�gS*��͂R��H�oi$�
O�_���~��rS���=�����#T�珥Or�˟C���
8䃝���۟g~�q��݃�g��Ucei]W��勍ֽyLF�v�ӽ���5�zsO��4̴P��=�H��Y�E�=*�(&HD�F7o2�@�s'os�ya�\�*y}F���v(�їb��B� ��ly��y0������W�?D�H�ob:g\z�S�>�������ҍ�z>gJ�i�l��]r�4���Eu&7ǋd����������_N�r�D�//Z^�UH�!x�P@��4�H�/!�'�&�/%�7f����'��#�_r�3�~���_W�����x��z�-�O����gm�U�ZV�Ǉz:����}y���}/��_�fg��{j���b�\,V���df��=G�d��~� �O�2&p������� �jG�~G������� ~�νk�s'[�?y4}6o���\�d6���=|�K���g�%2���ZЀF?u^K1 }ٻ���-�� s� ^}��P;@�q��x�{��+WƘ!��3U (�gv'e�N��v?�o�W5�'�e_������������7g<������皦|�q�L�4�����껓���� k�ɭ�3�,��y�~��gȰ�<��?ߞ�Z:6F��I�[��L�浭9"�����G����>�f'2*)���s� NNT�H�P������ϯ�et������ N��!����ݲ�=�9�Kы �}�����>}W@��4�)I"�;O
A����G�ό���	8��F<����?��9�1�g��;S���6����+��eS����f �llO-���JQтK=�M���
=p9�~� ���KMm�019��������?��چn��eF��|�S.�(e��X��[ɻZK"6b� ��N;�`֝��n8Q��5#�x���� <�6��ƽ�H� r叡���ݞ���GQv�}��f��=-�iGO����^Fq:D�6s��:ٓ��6`e���`ȷ��&g��1:�jM.zqǨ�Ǿp���9r3D�!�R�nX�c{��ڐ%�R�E*w$.��Y��/���+��]@��������t7l� �i��fv�w�}qumS���Y=S�]��r#�l~��qճ�ݱ�5����0��;a�4�g�wY�k�c�F姤�J�G�,��Q��$z>��� �k�#
��Nw�`IV�Nr3��]ǬiWں�z�Yc��'���2ȳ�����
�]��\W:��;N�<{}�>�{��w�^��N�{��##�;5�`g�ϰ3�ӝ-�jη�ꙝAY�k4��<����vv����1%�l��wP�$w����å�sY�Z.��-VI�CV��a�Ww���_'�Z��2;H<�	���ӷ���w����������OR�I'{����Y�*!7g��Ƴ�ĉ�{�����謯g�;�7����WW�;�]���-��yz�'���B��5-/��W���C#Pֺ7�+�jԎ6�����޻,�mC@���zK�mu� w��U!�r��ӭX]�V�jr�4��ϏqЌ����1�ݶ$XmԘ�b�;�oUv=��zt��U�D�Xˢ�f{4�5�~�*i��_J����Vc�	j���S�=��d�����[�������Bi�a��ɺK�}��ϻ�o� ��B�7�΁�̧o�Syd�2��5��<&�UyG�� �sڹ_ft�J�M2�C>�7�K�#�^�q�l�>��f��D����zu�s�u��7_PuJ� ��2E�Z�
��lG^�^k�OԎ��Ў�� s��t΁�����c��=���z4�o�0���eh�ս�i����ҽ5�8����e��W�U��G'B�Z���Y�c�Z�˽:G�ײ4Kw��z5�i,�J�5HWu�%��q4�,'e���hhצ�x����l7C�S����4}ͯإ�X�v�i"��z-c���9�D�Q�ױje������F&k�szc�}��<G�3��o�_��~�}�-#���Oo4��徧��kt6���Y5�b�gV�4J>��3|�S�e>z��Πo��7ގ�A��q]���z���-/͋R­%F�G�X��*�*���*�/�ݑ��ٵ-E��>�j�U�E��#�^C�)�X�>ٗ��ީ���_��B;��[�ݟyu�,�jcd�ޕ��}?ԙ�T>\e�zOJ���Ԫ�D�2�Zwo]�~���j�Lt�VՃ�����3����>0��9��u��뮏����^`#Y���8#�H�Ό����đ����4ޱ���K�7t�N�j�%�s�����Z����d���ܮ��D�tܼ����f��9?�9Z�&Aw8�h���1�����#~2��ֽ�Z���v�m�>ic�Ge�AI%T��S�ݭ�� i[r��b`���F�7�� G5��i�֫��5�����-Y����z9mL��7l"�4G� r��{��e�_�wX{������{��z�F��OO�GGk���Kh�<����5=�#�r瓋��KM�����.�Y��v�v�}I�Z���b;�qt|E���{V�Qm���,cx�Wqo�ݫ�-��u�CN�^ͪQV��M� �UZBX�~hx�p�q%q�$rFі<�^�{���n�}ޟus�o����Ws:븺�D�q ���s��%��ptWI�_8�%���P��5tN�m}p��ۻrK��+r�j܅��ڢ��L�=@���������?^��z:��JeX<R��%�0$� �Oc�>�O� Il9���t0���﷌O�k�:@u���h�����z��4~�CDÿ��gA�0U�T��<�����q��J_�z�rG�_T��]�N�ڎ�b��JX����*
_!>3[�˙޲�*������D]�ӽ>��:Uիׁo���:�g����~ae���p��c�g��,��{����W�u?ԋF��I{�׺�O���t~���Z�su�SD[G��/�_7K��풺پ#%`�O��p����g_�:���ƣ�KWJ�4ϪJ�B(��ӄ`�m�{�F���	
"2sb�Ź��'d딴�Ee��1���'�����Y��5q�����Ϗ8���~��^��t�3��Z�0z���-{�5ކԱ�-����]M��P�^lq�4���a�r���tHoOP����ab�M�t����F)<qJS��.֌Ek��`h���O�4��ݝH�R��[�+k�S�N��'� ���n���y����@� �ho�3�s��Z_o�4�S��ذ4,���Ojs�*��Jei�������酏�|�V����e���f	�ϟZ�𷺷��7f������fP�G���A�� �Ƈ��}���ۻOKڛz��ڔSL�t�Uc���$��y���4���i	2��F�v��7p;��~������t�1���^��Yd��/Oet� N�a��P�VN�7��FYZfu��<�<�!�2)��|�\�d�Y"������(Y	f@C3�Fb���r�/
،D�Ft`�ݞ�7rn��
�$�`r���1��O��[�{3���\Y�N���~P�}���0N/Ri�����oԗ���K�����v���|�:��JXꉚ��L{���YӟA�B�e�x���2��D���1'��/<����8���쏷�r�s���Po�vϖ������ ��xc����S�Mc�����Y��3���vW�V�r}| �7�rI� ~��=� p��,��g����>�ᝆ���}��m�^��Γ� V�ܾ���{��gM�?Ukf��a�S�v�P[`v��%�ge52h�e��]�L9ʴ]>��V�K-:H���l�AR��q����,z��ִ���"��>�	c��#�?l���WD���Y��>ORcf�'��[Y�Yְ��:�f!�5���_Go'�7|�d՚x��J�ͧ3խ0���Β0	���r�n@�n���m��4�q��T��YH��w�� Fs[�	쫰�����Z�u;�r5һE�֙��g�?�e�_^�mg1�R����t�j7��k�yK�'�JwI�Efs�=�߼�a�N���{��y�E�卖(��5.�p����"2;U��H�O� ���Y�w;���KQ�:����X�hZ�'A��JI��DT!�Y'.D��glֹ�w�)ʵ�BT9fn����� ���y�2��]�g��!���*8�� 3ϣ�f#��t�����%=1��-0���G��5���x���;|}U蚦�v�U�D�W�Hi�A���o��O���Y��/�����}�'�����:!�8��M�7w�L�\���L�VQ�O��Kc,�V"���D�1]���Mw5�~I�����*��v�b�{�f,.�[U��f�D��<��5$(�S�B���s�M���Ǳǔ1���"5��*����9P���X'�6W�%<�~b@��kU{]�j��%&��7�wa��m� }1����r^�)�/,yƞM���[���{�c��s���(��$l�m8�l �����|����CʍUEo�ꠅtS�c&cQ��FV2ȳ#���XI<J���!*f�lF��0�s* �E�ǳoJ��N 3�j���ݼd��dY�Ѽk���
�yPx�sKK��ia��~�;0�Ǚ��,����r�eG��jD�9�U[�6(�La/�l����bp���F��^I����̱��x��_匓�*�e�5g+f1tC8�=���PD8����y�%Ǧ07ǧ��F�Ԛ��J+Nb^f�̻uY�]���eV2*b���q�d$K�x�N�� ��E��3�,^�r2�2N�T�	��mUp%���Ws��
��x�2���lO�1�\�u��ǒ�� a���2HU8���fUĳ��b7�5����j��mD�Џ�I)�@�xՙyq� f2\�٦2�ل���yH���
�h����M�M�b#y�|�O���9�O!�e��7���i�r\�J3�Y�T�ݘ�J��6r�ފd��D��6���#�m�c#Bn#˒���*����2?mQf������ /N;! zc�E��fn��Y���)�8�`�����+zc.^=����.�;Q͋j�M&����%���f��V07VɐW�w��PZH��fՍbf8�����2Q�r������C�g"+[qb\=DQ+W�$]b�d]��D�+�݌��"Ś�Y2`�5�vɣ#�5�&�B����׊1�&�4��1ʅQ'�yyV^Jm�-�d��H@X�w!ر�!Qլ��zME�yZ�>J�'Ĝ��ͺfp�}1���/�F��챴�qY7	�X�Gݩ�,�H>�/�1�f������"э�V��Wl��ɘW�ߒ���Ȱ�1���<��vd����5^.�+!�V���ʪ��כ|�����m�Q��s�q�PfC��s��@ϸ
m�76e(�`�n�(��<U��vX�v6�XQ�f��b)�üռL�X��sIq_��q��q�3�q̿�A��S�I��.̄\��P�3�G9ּ�����ܜ�C���F7*1mF�錪�����(���20}�ٝ���0DTX�ӓ�&i��	Qb��� +^ ��<P�c�B�8H����+�#6�V�h�I��tJ��=1��n�/6f�WFs���`�㐥Z��$y82���W�z�49M�� w�J1�Y� �q6&Mǀ,K�Xɍ�m�FyFUEq�*�xi��\aPQ���}��^[��}1���)�;!���`l�!N�Z�f
�A m�S�i(�+��ExlZ����Ѫ�Y�/��q���Հ�m�&�悵��'ībΧ��C��a�n>/[0��~�2`{���(Q@���3�r�ݿl1��z��4�1�"aQ��Z*��l�Ʀ�Ă��U�Tm�M�o٪3"R���.��c(y�IT��A�ʺ��"#�SjY�hK�ݢ�)�3l���U�����EAa��$Ʈ>L�-N"|ýXBT���1��ܯ w>J(���H��2��P7�F�F�m@� ��ũ*�su��,�kQ�qʜ�b��'T��ɑ 3��(��d�|���Q�k+'7��fY
dx���و k��TK�$��7�&�:m:T�<��1ɦY��UI݌Ҍ�zF���̦,�1��6Td��A�O�����C�}1���c�۴䈪֕@�!���껇����#,b�x�-�U�>�%@Z�t4�CQ��s�O�=�� 1�O��)��6(T��[�"���@ƍ��D�T��h�X_p�j�H�$|��?"�,�J��u��Ne�`��eEM�����M��Fʢ��`��yNY7��Ǒe��^��Km��:4�*	�QȀ��8����/tz�d�l�>L� �,eY��z#�e�M(NAwF��?�6����1���Jճ@�8�4|��ݑ|�V
��"����1�T���1S@��7|ĉsP)��,ّU`Z�(A	cS&��aC�˲E�r%��A�@@V}���3f�Ō\�O�X�B�QZ�@�+0fwd&PUUo*5<�I�0�̫;ԩ>\�+�HI4�L�$Ȋ�Ee��7�rŷb��<R�P�y��Rc'/���tvDɷj���h���%��B�t��Jc�u$2����P�V((������"1��
�����~ f�)
]���wP�qC5b�\1�2���`i��2o�d�i�~6,��g�9�IƎ.-RͻrᏎ)kP7���蚶�hh�^����u^�X��ܓ�#��xǹ'��$���6�c[Ҵ
b��y(Uyg�-,�#��4�ؔ��Q�s�(}��v;�7~��U��}=��/�]E�8wPt�vz�;��Z�eeC�8]��s1�:}��\9�z��-i�7Mv�M+W��t�}��X���K�\��XF����Vl7p�DjN>�!@��ڎ�Խ�v��zggO��V7X�Gp�H�Z���:ǂDu�X����f�w�Y�=�tgd:��wc:o�zַ���Ӻ[W:oZhZ�j)������Н^4�j���m�2�f��^KC�Slu'���clj+�j�O�L�õ;��a�Q�-z��+}��bhd�J�)�>�}�����iZ����M��v���G�Qg�-�5��9;ge�c�+ Es�"�̙�=��������퇠����un륰�Ŝss:S��=�8�������� ��-V�V��a��xX�q�f�{�N�5՞�R�Z�� ���j_��J�yix\�,w�����LT��3�#�u��Z���l�f�ع�Z�"F��fH�E$-3�R%��r����D� �c{{���揤j>�}��o��w���Ⱥ�n;�ֺ�I���Κ��i=E��y02�zWQbe02�rq����Ɓa�e7\zO�kUwVί�têO�v}'��$�y�.i�<On���̵�g��	����n�m�"���:�������*��b��� v5;��?��1��aY�0;k�`���'������=G�������.���Yh���n�����}cS��ڞ�ɝ���.>��.6���e���'�ˍٵS����_ѷ���߷�I'��� �/�b�7s�*��F!GZx��+�;L3v����>��Ki��2Mm�h&��قɬ֧n��Q�=ۇ�$��b�L�bE��O�BvӺ��OC�[ُ�Սޯs>�ܱ�~��^�hR�n�+K�ul=G�3�:�A����ҵ=[�2�&vƜ�h�����C�.�R
J��쩣lݗ=mnQ�f{SU
k,)�^8旰1���"4A�"��|fU��؛mOt�8micx�u��m����l���$��X��kM#v#�l?����ϵ��^�{����p�g��=����߮[�:A5�BX�m'I�u]g/�z��2-+i��*��`^� ����[�=� �EsM�:���4鈧�麖�CZG��� ؞^�����I�*LH�˘�N��ײ4F��NƁ���oJ��^�4)�Om����c��ڭ�J_��T�ܯi��z��GK�#I�>�kO�.����]�8���c���5^�up�~:"S�:�Xi�g��y<�	��ΐ�]y�S�2o�#[u�s_Z�O��T�]�묖4˿.���O��b�'|��^���L��k�������5���#e�Z姺ajVL1ۮm,�G��j+��}�����;��m��d�۟t]���iC����������V���6�ۘ���e������5|�d䓓�c*���U��>��:1�4n�������v ��4��Dѭ%&U���cJ��J�,+�p1g⮇Ww����STٚ����V�g���\�V�䮏/ʹ�aE ����gg}��E�s�S��^��=3��3�]i؍g��N��{���H_�����=5�X�%�8��Zsb�ڮ>L_�V����w�m@��G��j�|�mXKr��yX��oQQ�`�b��U,zQ��5�j��hj���^�e�'�ح%�:Y�ud:�r��dKI�FA&F�^����N������ϫ&��.�{|���}����s�5f��퇽��'���֫������*c�S���_#K�K�:__���M�5-V��/���kD%�4�J��T�D5M#=���"��_��Nx�ΡA�}]6v�b����:�r�I$5�]K�a�x*�2�M2w���
�-�Q���/6z'�z�R���b�?�m�~�ڇ}������g^k=Oם����J���,̾��)��t��� �K���P��4�+�2iS�M��9ѭ��b;��/L�rCn�z�C���#����$�X�2~�D�"+�,NW�����Cu���ΧHl�y6&�����vC;�JH%��Ԍ)SVI@�&��^9#r���;U�"{}�v��Ӻ]sz�u����N�t�i8}���	�v6�����U��3�Ϝ�;�m�Q��;s�H�N��mA��OOӫL��&��i�����̨����4����ɷC��m��^����jvnB���S�{l�G�����N8�w~�Ĝ�=��q�I�[ڔt��{���������n���j��/�jmJ�t���5X�%�xU�W.�yG 6�C�~�|m�MC^��4ٶ&J��Ud5�	_�^���c��1*��h�y (�j����;���ӽe�ͭ��[T�[�Ul�6�Ij�N�G9�Z	���u�������Nj���h���o�����K�}����YZ\����������mp����v*�|�2h:��ލj���_t�Z��ֺ�����
�ԬmN�'�Զ%z��
꒕�Y�7/W:���K�lv֝���:u#c���e��շs�2���X�H���4��*ڬ�����JS�Z��ڍcG����^f����t�P麖0��;�4��v����3�]7l��3Y�ok�n�kX��rƳ�<���,�I<x�Ɏ�e{{�^�#nJ@H�C��KG�F�I�V1�HPG^0����������V�y��G�v�1�������K��9V�;��.��4�i�tCkqX���OO�s���z�RD```��LԔ���dS?}Y�)�<f�EJ�T���6�R$Gn;x�!^㐶������	]Hh�`\)Y�H�B��� �pI*���g��hz�B{H]_�'lE�:��_R�a����,�D����^=��T5c��J궙S��+���ښ3�|R��X��G���b��=z��y�bB���J���9� �9�~�����˷Zw~:S����z�z�#O�u{��:��-�ՙ�'��9�AL���P3ȴ*�u��ȔmZ�=��8��2�1R�������D���!pO֧�����.k2,������t�d,=+�����a�?Y}7����׾�-�y]ӽ=�t�E�C��{k.��,��!��P#��%5Jj�L�&͐������W"�d��nG5O���� ���rV,��o�He1J�AA:2��OZ��'�ձU��37��w�2���ywC�8R$H�y<��S�V����op���������@��'^hwҵMG7^��{�rtn�lx�7�J�ڮZc&�%��������6���=3��h�"Y���Q$L{��@���'�^�/�3��̲��1g<�P�����p�[��;�}q��|}�����A�ާ�.��^�����uF��8��p12f����M�� I�k��x�=�U��G7Q��Z;�lޝ��@g^( ?���$����s��9_N�T�h��廇?d� ʜ�U<s��3F1111k�1?ʞ(Q��k><Ts'�m�O���as3x� ��?�� ������� >� ��� ,����D(� ��3Q�,B6�� �_b���B�^Da�� ��������	��?�"�gQ{R���M�*� ���,����׍�&��^0��'���={����c�L��q�?OYh���Q������x�O�^�M���6�>��ja�f^���sϿ�� ��S�"Qǿ���� ��s$���k�n���i�o����\4"�Z>ŀ ��w>�2iU�VNd��py }�>������u	�? T=��O�����_គZ�����U��SN�Ȯ�a�5l܉��6S����� �r����˫j2�V!Ӵб��&F����K�����#��X�Y��S�� �v�� <��عn��h8�zF.723�|�]K���M�T��ѨGNj��P&���. @�ʗa��^2����<�(o\s��b�]�Vh&��v�,���a��� ��=�v�J�7�y]���/�]��׶�/w�n����jtF�����|o �RR��=+��N˭
�����OZ?Fliu}-���S?�@@W��W���~��
�)��FEڷPC��V�o�oݵ��5����v��,=K�
1�_���g>�;���׾~�}�{R��I��q��è;�ݮ��_��R`ꓶ���wCS��S� S��V��:�����&���L�7"��$��D�L�W�˚Ƶ�jUip��4k6Y�A�Bщ�ծb���i^K2H#bK,�Y�s�����vv�,U4]Z����N�Z�]�]*x�b���"C�� ��@9�������;�/�s���a��v���]��q�����5n����=��պ#7Q����t�>FF���S��2�jlf�8�|[u�p�?jk�f�����i7�J/�M^@Y9Do��$�+���FA=��6CS�b�U4�֞����h�U��Ez���ɂ��ϕA�� �zX��hv�ܮ�{������o�7�����_Qw�W��D�W�L�]{��TE���ޥȆ/���gb�1̧J��L�/Z����3�Λt��`u�pm3�� [y�v���Ÿj�M)?bj5�M���D�MJ	8|p���v�-��M���OM���k���̮�zKIb����Q���kR,�IgO�,�jeK9��K��@��܇@�E�rs��S鎔����=�?A��kt�O+G�\\މ�S�=#X}����l��_�.oSWM��M>��U�L���� �ޒ��D�vj	��Zg�4P�r���#�.�SO��mI�7i��?�c���Eٷ7����ܖ}RX���E�="�J>U�R�ۙ�9���٣��� ۗw�Џm�c�;h���_wCV�?+;/�����·Q�X�n�uө�i=@�ն�}O;+	'�ZR�,��������u&����T�DQ�n4�0 F4�Q)���2Ai�U*Ñ�qw7�� Lhi6�揥],�K,�RO�n;�7�V��0?���y$fp}}��0}�w�۟��r�s�=��f�Ԓ���4~�ѺkZ�M.z��Ӻ֍Ԛfn-u�*Rs|�Ic���VL��u�;kh�Kt�k�^���N�w0��6^�B֢�)�;(Ѵrf��Y�Y���9)��_qt~kZJ�m������́/�<�h#2�H����CD�0+�zoaz�������n����o����K�uV�۝�:���o�z\1��t^����&��[I�2-���f� LLJ͒�׬Z%�t�r[�n֫�5�Ւ��a_���3y'��䔪�$�������[wK�D�a�fۣ�~Ϋ�Dl��ܑ��]��xyHA���,x� �%
w����~����4m�ߥmtN���s.��zN���1�O�]���e�'ֵ�6��t}YGMº����ٟ1�o_������}cr���j=I�!~f�"� os�#�wfc�X��'�:�I�=�m�+V�41�c*�����P������W�1�bH'5��?v�on>�;�گk���ChW��25N�����������/�]�A����E��Y�Z� ���ZE����ޅ>��&���M��Y�{1�]j��#���rȞZRM���@���Y���z˫����GF��Zz�Z��F�h��#�!x`�CcƂ)|S��4�!4*���}�h��?}��O~]u�w��'ZN����j�M��T{�E�~�����'+�k�2��5�\\K��i\زQ�Wt��I�i�Ҡۺ�&�]1k�nJ �ͽIjw|)R�Ww�`���,�36m�Sn��Y�l�m:׳��-^+����[�k(*�P�<�2�!�N�����I���%�ٮ�����u�iwȶ��W�����K�^���[�����T�ΦM9�T�N��\g�Ț�؍:��z����ϑ����;G9|�H� w�9���t·&�Y��NF����������9�J�>]T����"T��0��5� Q~����s�������OOtޟ�=_�ޠ��-G�=o�L�}w��=�N�i�k_��>����[����b]�ъZ�Uu�6í�2U]ah��Q��hO��N��!����@b,�)
x�����;Z?Lt�ܖ�J�\��LM^�y��;���a?0gi)�?��#�3���+׾�r�ý]�u�����j�hu"fh�};�\'��n�MGR��/�`Ůɉ��z�
+a��NB@�d��}堾���J�M�hvޚ%+5���DH�?���"�i�C�/l}�ӧH��l�jۼ�A�7dIR9=z�����,�NHG�B�1$�$^u�n�꾣�]w�z�U�zi����麆'o�����{N����q׶L�l^��U���+�5�O��]x�gJ���F�F�A�Xp��LDoj絁���;z-BĮ�#8�X8`9 �y!�v���(	���7۷��Λ�F���u���즿��ףun����3�������{G%�N�`��g��4m.n&u<�nj��U(����h��P����1���0�Ї�{����R�����C��G,?�	��,=g������.���^�v�B����;[mE�;۔�L��k�9f�}M�o�^�׉x.�:�1<]7�U,���9'��Kz�q����<��9u�,Ǔ���� ��?N>ٗ;a���%���������=YM:�ނͧw����)����8����⯑|�mN��><ٕ���Xu�9��������s�I<HX)!?�?�<��}�3�]��_O�����;۾��ޒ�v'O�?ez+3��3�un���m��O&��fF6��f��Ȗg�#<yq�D�2��q,^.����,��H!�d'��zv
�8n����~]E��:�1X���#ȯ�#�<( �A��z�����=��F�N��:���{G�P����z����q���t�;�=��|_�c�˪d��#�� [&��بV�c�N\��ۃ�C�(��F�p�8ʽ:��s"�VX��][���B9��@�P9Ϸ��:�Bv�_�^.v,�q{�׺��������,�� rm���ń0��=�{b�S�3�Ŧ-��B�H��fgrB1">�%�b��y��<���B����������Ϣ��q�q�x�Eg	Nz>�;X�J�- J�?�W�[�*���}� �c�qk�@���I�
��$~y<���q�//�im��w�x=� ��<q��Ny̮��t*��)�ɜ�ˌ��[�EQ.,��
��~�޳J�wGՠ��@�ґ��J��^�^8�� <�lj����2'������߯����6���j�`k:`�<���H��8�rG��KJ��>�v�.�I���J�^��ipv�#q��i>��p>�����U�,kR�{�sc�����_�N~�흖����?����#������蜽3�����uTkQ��F���N���5�KE����ujZ�1!���4�Ni�%�M_Q���~j����:V�N�_���9��{�H��[=�$2������
�s#��� �?��_�:v���o�Cմ�R�Ϝ�kP5u]>H�x��k-:L��a�O'�a�?t��k}���Ivۧ�ޫ�����c�=�Һ�+����h�L��������u~��t}W#I���⦚������t� �][�:.��6���!�fk�ET��M������{t�S�7�V��(�\|��$�տ��3�Z���7r]�ִ(V��t�٨�~/� E[�.C(x�-�D"-j3,�O��ަ���Lޛ�]K 4�.�z��>-k�dc�ӭk��ݼ�f��]�Kr�Vmuh�4=N�s�P��C �)�?ْt?�>�n������J�[�Z�}wM��|�F�s�횼�qOn>�����fsi���h�U.$���,�x(#�<A�y�l9��w2\��r!vV�7t���
[�زL����9rc���4ҙ��.N;�dHrq�1q�Mi/�d_��(�%]~�C,zcQn��;�E��,5 P)Tb
�^m�k9v����*�1�����̆�,�� ?��7j�E;�0-*-�ʨq�=R�|�P�'Br
�R���H�0�X1��a���b��h^�wL��?�J���չpRK2䀯�1լ�|i%��4y�-$3D��x��K<��3qN~N m���6���DJ��ɌCO��C�!Ϳp̟�ə'c�,c�Tum�N�ߗ���4d�w���m�!y)%Czc�T��^=,��O��2�T�+I�^hSa�b�l�LǏ�9�8����>D�#�8���#�쪡�u��b��,��/qIs���4��xm^cdQ�B���HbʶLl��c���`p��j��dVs��},ł�K��2�,c�f���m:9�Z2D$�2m UQWd<9��zc���IF�lu����艏ǚQ8�+>^?��@B��K�5HHq�:���p���i�F@4/��ܹ1���3��͖y���E�v�mT0^���&N�7%X� IA�T��dO&K���U�"�Vhj�[�P���~�c%6�g�*����ڔ�����H�ՊM�q<��1�&�ċBx�I�y�-:F؏ʎ��.EQ�@ T�Ȉ9��[$]W��h��^Bk�[��5�A�>-�ʒ�  1��ƍd�_E
㜄f!�x�i�\Q�2N���I�Ȓ��7r�E�L[2c���L�Rr�2Ӊ�Vd  �_Lc��o:*Y�d���gvUƓ�<ם9���J�o�T�t�K��d���։�!]]�32��gɳ`̬c@c㣎S�$�CQ���Gv>9�+�<�Lcd<�^�3������6//�n(TI�����ȭ+�c+E��+E��qx+d;�L��
�/��G�D��4�C�B�bK�cpc*	X _-H�+g!_�Ք"�=1���Y��Ygl�ҙ.�1�dqO������`c*�^���%'JU�$�ΔR��ݹ�c�0�#�,���/o%�V��$'Tj�)����0� �(r����EFX���P�.�.�HJ��PU�
��1�x*r�1I�7����&��%�Ɯ���v�G�Q)�yUKp���l������?=�����Ͷ惈ٌ:^�DUV,�NEN.<�Q8;ȰA� qe ��8X���B&�V+G�$�O��G*��K�Y���.D�r(9l��M�̙�s���� oz*�?a&dEB=�D��"��$����#�>{r����`X����d��|�R��~30��̓�7!��X��9d����Ӕ�A'V\���7!�{�˹���˺R���N���!]/! BQI}��(�x�eFŌT�T[#���^H���.D���ٛd<@$�v�pX�J^�x��mgy����M� )�
��y�m��Fۘs��2i� �6��炅�d��99�6� �@?��~-�����/Vd����(�S�"���QV`n}1�7 [ɉWW��g�ݩnW��)� ���^`E?c��W���T�ɣㄢwD����h��7+d��c*I�YBJ��x��.��(�!J�?�&�&��d��e�aX���̷P+H�e�H(*�y�
�����[��1�̴�lx��(���&l���^,��ǻ���P��l?�Y� �y��W�Ķ}����Wt�������dB���*T�\������-S�:�W���v,v,b�<2�\��>AwJy#"M������dP�%p8�P+��(�'ٗ!�(�W�5���<�|�YI}��c�����EY�a��� Il5��
��DZ�0n,b��d�Q[�c\����G��qέpT��ًn�l�9p��&�6��ᨛbN�4��}:��WĜZ�J���lw��5<)�8����1��_hC��\�#Ƕӣ���OLb>J�f��e�b��sV��*MAf�W��bU��ȹck(���9�{-9P���)0�L��Ls��*�wNLd����;cB�\P�[x��[YmE�7d3W��7$��V1���m<zS$��Sώs�^,�gJ�MD�m���C�Q��V3u�stn�+��R�P�&�cH��=k�dJ_�O�#�xW��"H��b�5�㻺�-}Zڶ��}�Z�џ%���M:��H/�h����ǚ�ֿ����h�h���@��x��^U�)�� ��T�ԃ� V���ץ�3���{�ߜk�]��uOF����u�b�V���Y�Li
F�-��6u�f�w����A:#�t�����{m�,̭>�k�{W�m����8H�CFX�����i��C�ϭiT~f1�������h�y�M��yX�,��3�x���ՠw㫿V��~�鞤�����3�Ρ�� ^^��Ldt�
�U���迎�,x�ZhQ�O�� ?�~��wp.��I�H��-��T��c9�Ɲ���7l��
�b5@��������=&ޏY��;��X����u�CQ�@"Rp�b��t�:��׼?u=K�3�$��%�]@��}�����}�M�2s���uI���)���a6�3�a$\�l�d�M����t���z�,{�sܳcS��'�H6�1
Cp�QT�$j��T��|r��?9n�՞��F�R:�퍻�V�J�S�~^-W��i��O%�|�4kאD�����=��G����x:C�'Ytj{'�jaj]7՝K�~���Ok}�~���ru�;?/���e<Ș��퇑�ke-��:��n��{�[Spj�k]hlЫ��]�)��"�h%�Z���x��K1,ELۦ���z_T����m-�	�P��<��\�z�X�V�QͦξPE��A��S��y��_ڧ�.���� �n�{��9�ٺ�pr�������N��\�[\MQq:�q�p�:S�"��kly�$I�i�J~���������[u��l,�sb�mR9C0]G�ד�#z�f��o��s�n����.گ��=���#�:�lб�D^�E]���[D��x f�{��׋��:�wf����:�LN�������.��t��3��t�Ou>^6g^�nV���	���֮c%`�������tOE�zkԽ�[T�5{sKf���Nqƽ��Ef(�Ĩ��`,F�_�����4����.�o;Z~��VH�����\Q�I���b�̲J�W��<d�9�:/�:�z�F�����Z�����p}�{j���:���a����ܗipr2���,Z�A���4�Hd�
t�3��uo�=5���u���?�Яޯ~��ZQf�MV2�DP���L]�N�s ������;���w6̊I_]�Fm>�S����Tӿy��^g-b��`U2Cq,��_|~ֿO���#�]��W�ξ��s��7�Z6��޻�P�^�/Vu�ڮh��/���y� ��mh�	V���6``Δ�
��;�Z�WP�����&ҵHlA��Es)SWY,�R1>D��ㅚ`@c2u�v��ٕ.˵�nQ�����,��*��.�ߎ����;�T$���u�j��ޮn������L{�t�v�ێ���v������O#Pm�t�*��yڸ͎�vϚP�Z鋋�����]l�o�^ٗ������2�kX�u�j�ݹfHZ�,�VX��cFH�(lXie ���?Q~3����� U��h�WM�y운�JL�y^�Q� �<�[wR�+-z�#F=d�OWv��:N�[�{��}���`eGT�����>�;Q��E�M_I�>�:D�k�E��ei�����V����%ai=H���m�;&�;CO߶"��*ݖƁn��9+$��Ɠ����/��D�cG�*��W�z� KWM�wՋ��ǆ�ʶ���UjG�l��k�]N���%�d�J���,�����;iԸ��4����=3�Z�_S˽���P���uN��2#��6���kN�թ�U����8��|�Vv�]��Ǳ�	�.��$ۚ�걲wIC����!�#�#m=���Î���'d0�����'{�{)5�����m/���TЉk��c1��;Jd��9�&�z�¿9�~�pO?r��;e�{܎gt:K�u��/G�N���|�+�=k}]� �����h�5�;U��*����\ŝ�l���ֽ��}�j�RƯ[�mN�=$�ކ{Ms|ʔLg��C#3�Q2�(���@�.���д=n
İ�K�%g�Z+л�K	�-����+�'�!!G'�{h�׵���Z�W���w{���4��4����ؾ��=��?VL��Ϻ��t��tҴ�k�-f������-�*+���5�궖�56��=}>�Q�=J��nD5j�BI+ى�(�v����<O,����D-�G����Q۱ٿ��v�w��y�L�Ȗh�!�b�]k�I�˪��=�v/T���w������>>����u�o���]��4H�Ի�٭c�o��X�W�VV1+:�-��v����M��5	����{#w���EJ�z�=Y^r�M6d�:�Y���Y���,e��3�~":��v�8�G���[Q�kXMB�:ΐ� �.�+I
��&�����b1��Op��{�w+�>�:�[�\��7���+�s�����v�5�[�z;!�'D��
��8���Ȧ��֩�^������6F�/�v\�\�`�,�'1�v�RY�d��đ��>�H�*��/m�:��_	�7��q�ȱ�R���ѫ��u�g��͢X�ay
4Ͽ>ҵ���Ov���w/C��ڌu�u>V����W#;N����d�R�)��_��R
��3/Q]���BX�Z��!:��/d����-�b�d'�^�9%h�U��Mᑸ��ᕑ�L��/�{��s�'�yA��:/a�?�^�����{���i�����:�3O��ZZgNj���?Mc�t�4�@À�.#��'Oŷ{�ծ�K�sb��$�;JH}��v#��`���ω4��D���C(<���@'��x<���^�{��/p]H5n�ײ-�h�x�_E���oE�F�8c���leVzsX�k�Jd�_����I4��ؕ��C˻Ic�'����x���*�(�U�G� �{��ǾI9�]N\.4�����;���o�  � �~��ܣ���h�������~���� ��\��eB�L,�ًQv�q?������D� ��9� �� �<{ϋ'���?��f��3�N��Ѻ�u�o���E�SG�?/J�031�p�O�0�5��b���d�K#N��}��s恻Y�Y~ݮ��to`��+}��YH�#Aj1,=܏_f����U��]e<A ������W�t���Xgk�Z?Kh]?�Z*����DizNf�}ӘІM`�X�fZa�O��s�z����gvH�����} NyD��Ԅ@O� q�<�a`��9w�?��=o�.�f���Y���K��ة;���*���m� �v�S����}�� ����ݟOߏ_��SPS�G�"w��#qB����� k��ײ������O�s��~��҆�BG��� <�k���$թ�~w�Ыf�ހ���#��+ĥWȿ�=�9� �� _g=Mx���?r>�����t���mO�4�>f+Ƶ�}��@8�E���ŧ��m����@���Q�lJ�9�<z�x �<���#(Y����x��s���?���=�7Oi�:WW�1n^��1t�)c��%�u,��x�����,��Ӛ�j$�E�L� }>��~��?�}`�<�n�9��� ����{�=��d�h:ìm��d�ɲfօ^l�4��pE��T9�l��	8�n-g���E��`�y?f���9�e�t�
#HS�O?sǮ����x��Rbt�N&��&��*Fjo�z֝�Ԝ,�3f�
H,o2����8ںz�"�T$��Op2�N�ѩ��?�� y�oZ2�h��K �1��oa��� ;�U��Y�9>�;٥��}�vw7���}��i�mwV�4N������M�<_p^ڟU�_F���.!��b�]+�6�z;~8�߶z!��7_��u"���3��o1�L����Z�Et��
�%�HĨR}�{?R��SN�&ړ�baj���G� ���X�W�%�r�u^�]{�����J���|^�=�tf��wk��G��'�_�ޡ��_B�Τ}7Z��zǫ�=[XȽuܥӲ� ;*Pɰ���y6�N��T�%7�Hw���Mu	*i[ZܱZ�X/Zp���r��i���ps���ʾ�S$���v�U�Ə������\-V��,3,I%��i����J�,W���y���=�v����uo~�)���uc=������g����'�'��&���������=�i~��$��2�-V�m?U�9���.�[�����~�ѭoQߑX��CO���$�f(��9���s�IYEf�	46S�����A�-���Z�T��Z�iV-MkN�9fI%�R敩)����KLh{������+=��;u����j��Fv�/n:3�&֘dW5�=b���{{�ER5�W���J��lg4�H3�g�ε�m���*�����X��\�>ш2�3�I�'�T�K3�%��� �n~���;F�5MǾ��7[Ghtyt�K��RB�[j1WM飂W��X~a�_�7ݗkz[�b}��3�?~��Zu��vcE�������J����uw3�q����ެ��ek}E*�j���3X��\:���#��[��gR��Yہ)���^���$5�Z�d�H�i�f_�ӨxS啧�i��{��5۝m����~*��Pi�5�چ	>fx?}���X9�z�� ���B����}����?;��׳����gt}�kFI�oz������R��F˶M&��i��چ���yzm+��R�ɤ�F��ćS�~�ж�/Q6~�.�v��+�B�	v���<��)3�a3bxp�"ωχ��m=��n��ɶ�.٪��^��A��/jV�����9�D�H�4}��L�S� �O�tV�m3�7_;gc��zV��z/q3$��#��?�����n	��I�΍�=����j����.d��La'�IxZc	OC�e(8��I~#�̵��5�|�$G���Ac�9�"��$?�̮���0'���czOH����^�=�{a��x]���T�b����X����n�얣!����Иx�z���T�jD��\���_ǝ�X�W㓭}^ٻ����iZӶ~��:��A��t�Zi#�c�fI|rH�+Vh,ô�g௥}+�{Tnmѩ׳���KS�hd�-���&��-��v��G@���?/�.i�Y�{��;}�{�����~��붣������+��:�
�i�v�Z�j�~6,��
f6N���\*do��R���w�Ԥ��V�Y��/Q�E�p-�� N��0H$�Dc�>)zu��hny��N��u�Qؒ*���E���i�
��	�"�	����9-���Wyz"Zm�����%��M��_V�G���ST���;�kIr`Qt��Ɏb�X�X�)��u ��m�Y��3A����T�Gf3�귧 A'���e'�jЎNr�-�������7HxL7vZ�<�-�/h�+2p�-���3�^����v�������>{a��[���M'�w��@n�tvu=n�鉦u��!3����DN&}�3�MY9��Ṻ�Ow�ە&Զs:{TO��h-hʽ�L�%�$6�$�V����^�|h})�k�n���,�G�Z;��G�~f:� (Rj�ܑJKs(��>� P�縭_�G�~�������v����l�ס������*��ӺsU�� �]G�uI�kQ���������%e&��O�N�U5��i��(�MF��DrWYt��֥�
�g�wm� �̨`
�$|RGҍe�V�c�Dӭ/qe�.����i����k	�Yef���t��ϼzt�g[��d㉤`kz΅��u֣����*���ӽ#���t�޿�%9�s���V�u�>�t� ��M+.��w��
ʕ��}&��pІ㹦]q���1zu����(`�N��6� ^�k+���ui���9RH0�����W�_{>�;�������i=M�>���gw��K���#,&>�՝)��"��a����A8�ŀ4R1-�M�u~�n�[�x܍� H�/rW�
� A�x��,�r�V%�voC��ch]5�1m͡U���d���ͩ��ԡW��>(�����3�������-��Q������ڞ�?F�����6G�΃�.��Z�Eu��ˮ���Ν?+#W�3a�*x��y+؝�$�&fXvE���Aʎ��*���� �s"+/��x��r�+�VF^�9`G,��Ͼ��G�lz�w����=��o�~��]4��/��Cu�e�=K����t�V&����13�Dĕq��:�1��M|Bxi����x��~�)��rb�;�����H�м��ܣ�;�fW��������Ct�I{��A{��g��N��^Q�z����m3����33q��2�]/������pt�iB,���FR��yb�;S�����'�?�� �>�ܓ����� s� �u㱽��/���tMh�V���p����>���R�h�Д�}H~���C�����2+<������Jlș.���j�0܍ɞAD*!�=Ź��9O���~��^y+�����'������܏��w�z�l�;�܎��c��ZZw#�4��u]u��ޟ��>���gL|�g�*XOZ��D7T��,�	�4;f|`��f�Fh��Sq�1�{\v�\�i�>i��4��!#��Ub��F}H��Ϯ�|f�:����G����u�[u������GH���u&?�����p򺇻X���{o�'U�,_�Z���1cO,,�SW�ϒ+�ĎT�e�W���}px�>����qZJ��a[�� �؟�C�I��x?��0�t���]����λI��zm��	�b���}��ţ���>r����=�n����ެz��{�3�7�Fq���1�l���� �  }�R����;}�#���q�'��k?C=K��L,�6D�q�ı�V�m&$�қ�؅�U�F�.�h�:���l�Q�}k����{��=�کRz�h%����C�� ��y��/[��VZz�0Ɋ�#�,K��� F��`I�ߥ�Z:��S� ��������O��e�7��YJ��;���O�?���Mq�[ڎ�=k3+ �W+"��7��fE�$��������j��5Z��z��Uy�~����fQ_O���=����/qfb�俓���.V��g�Z���p=��[���ǘ�"�+�����oW}��رz�Q�i�o�H�A��?�@��y�n�B(��f�����O*O�� �{�c�}gD?Kv}_���w;;��-o�WZv_U��^����G��9�[Қ�n���K:�v��՛F�tl�d����IWp~�Y��ۧT���ޱ[yڴw�D3*� ��bCY&>n[ځS���4� ����n�՛V�]f��*���ԣ�g�9�-UK2W�5/{4�b��Ud~��N��;�4����ֽ�t޼ᴩ����g겈gMS�������r-�:ɶU�(�r�1K��G6���cpo�BĄj�Ԉ��-��ЅR�"@��*��F�Y���F5=�Ӎ&HԢ���Ә���~�9׀;gid27�3��.[���9����>���h�Ӭ�I��i�I�ٚN1h���]��}��q�Վj�RD�%�<�16��o�2ŤޏPۖ�%j��GQ��deR�ŻV�1f
�~��ベF��?�n�K>���~�8-l����і���ϵjP�
��΋�a$�:��~�:sZ�0��6�̹dANtM��g$|pE�C��u�ݷ���� ���|n��,j�?���F�j���
�M�h�EuU@���c�1͔�_�n��oWE�=d���݈�a�J��(B���ŉ�yk���t���+c�O�~\+:�y��l�8�bҊg�M�*"f掅��Y@)�C-y��b&��v)$r+$���$F���*�0?p3t��0�f��b������Õx�B���ں1R=�q^O��1��,�Tc�Yq�М:b�b����מz����r�b�S��!�������x�!vb�G.�X�*�1�.Eԣ�rU�(�#s��'�Yó��6I�2��q/�3H�Y�<]�8ʯ�d�7Wz����L��x�Lc�$.�KH���J65,��o��*�[��8 ~Bn+�c�r$��1�'�>2�@�mۛ5�����%J���?�rƘ�Q���5L�$��������!��b�ao#y��O��VCȎy}�� O�0`���l����8jі��Ev�a�1ww_��.�n�x,aQ��Q�ޖ�o"�/�]ꕓ;lT��oɷʖ0��Y���᧴��V(���!�M[�3��1��c��9b�+,��&&[e�J�vUf�����LbQ��i���jj,1j�\��u���W$��frޘǧ���ET�V�U,�Q�D�I �F��~���X�73�|ȋ�,��`<�^Gb��Oi�9��c"M�D��4��^-�+V�	~D���Bс8vR7@G�0�B��R��T��:~D�@3"�c��y�[.�rx�c&�So�ԩ��!�����'�<�%�ހ��]>����Y}1���.iifdE�ӑ{.��ϖ;K��Rp㈧!�Q���vc*�,��ڃ�X˖$�8-Ğ{��e^�������T����:)��RW��[7���
�/	��JqP�E����[<���R�.B��b�s3e;2��%�2��2cȳE�KH-E'Z�m��.�[��$3,ׁD!"�c#I���3�$����N
'
_��LbE�Ҫ��i4cu�7�Jaf91�w�n_�E��F�|��Ю�`�0Ȥ�Z�q��	�i��a��*=1�e�P��]qN��U2O(sZ�]���U�_,��1��d�7��L�ڀh��b�d�'5eN<�X�*2�VO�L�7���[
�n(�\,����7����B3�E����ı�NkG�dd�L�+!�Io���B��2��)b�)2N�4pȿ�o�,wo�bө!C�7�����7��c-␎T`��m<w1���x���ECM�EP��)c���̳� _�R3�q��]ߓ,�t.�o�2�Ld�d��9~G��$�Y�u�K����Vr�͟��@O�1���FE�'�����!YA�'�8!�AI>۫>����nZ�uwC�QK7� �`<,�,]ڟ^ m� Q���7^)=�/c9����Z�x �ǚ��E
� ec�1���9X��P���1����%]J�RS�
��W�S!	w"�fQ�-4���>��ݕ[�|M�,a�����!��Zy� 7�ҭ�q�ANJ91�l��%kL8ZOJ��(�D��I ����+����Ō!f����i=|Q�D�]l�Di�b� � (c�ZL �I)yE�������Ǒv�[� y�ܯ�2l�B?� QH���Kc?�N�m�Ǧ3ΞkUՑ�f_�z��U�PK��� ��A������H���5r6�%�@���'��3U Ú�8�P�cp��d�(e�%ǤU9y@�d`�6no�<�m�1��P[lh�y���s�ࣜ]՘�O�Q��y�Klch�%1�.O�L�8�c���Ĕdzdeb���~�ܖ0X�H�iP\����N�����]��p7�N��c%��H�3U�5i<�V��W`��Y�$��8��b�-�;Cx3��E�$���|�,�Cή��Հ�M�J\wܩc��)����S�6FD�#���Ha�TR ��r>�Ül{�~^1\��8�%��k<���>/��f����� L`eKdAح���@�*�����3̰�]�f�滍��V�HV�-t�=ӕZ��Ipf��R<�=�L X��<�*���d3�M�8"c�Į$��͎x�t��6+�cԫ���^���A�(�^J�w�Q���	~nG �L�O4jY��fDǺ�J�72�mlv�撧M]����
�ZY��)�F���yZ�>N�>6ض��+�m���IƣfpB#TK'1�y2ʎA�#�)��� �v�N?c���ʈ���  I$�  {$� �$�>]���" ,��UPIf'�P$�@O��c�Ƕ~�{��sB�����tNV>�ם����ܩ?.��M.�_��r0�;�LK��Z��t�`�<�wukM;é:�~}7l�N��M���hX��B&�����M0��[��r�3����:МA��`�����Z`�fUsc$�'�xD�M�ջ1�/{N��>���'xr:Yr�z��_�u�ۮ�հrPҵ��s�~����T��C���r��Feb������>�y�軪-
��$-��Ogb[�ei�»��ʠ<dٴ>�s��K���}~�Y�k7��J\w�Z�/Q+�]^h�X{;pNw����G���N��I�]{M�݇��힩�k=UКֻ��6�bixz���iz����c��3[$�,˂ -@ҿ��k�g�V��R���nYF�ij�`qa#��#��r1Q�	�P�PR|n�Αj�m瓧�R��	%�6ň%���܉]��i`��G�?P� ao�[�4|�c�o��mF���y�76���6�ӽI�J��]A�
c�y1�Th-"�<e�΁��J�N�w���ۧFX�ځ��4rw�Uv�	2�~$��c����������j�n��_X���:յ U����h(��0x��� b�����Oh~���v_�7x���{B���a��S�u���q�N��OҵmcLЙ�Ӫ�a��y���!�dO'y��7����O��7n��N��_�j�Uo/}�zY��WbՄM+4�����#�ٽ_�=5�>�Ӷ��җN��j�J;%%+<0�$�b��a���`J>~�O$�$�fCڡ��[vϣ������g����o�>��z���>�^�����|��Ρ�i�o�(i��ʻ�!�2�3)b5o@~�Beo�j��m���.�c2�lMmUc�V�xd����2f=Ѥ@1tʺ��S���ol���m�wN�>�H�( �:�mY�b�pB��,Q�w�vvɶ^�=�w���b�ҽ�{��k���2}�w��l��v�S��'l;��M��gTJ*�	qm�X��oW���эջ��vMKf��.��]�=l��=ߴ4�8[(��껬�8y 	��N��ô6���N�Cu��P�C���+��ѯ�KQh��2��oM�-k)���w��o�.��n���u �F^_�]BC��Go��5~� ��ؙغEz���l���ҵ:&���-3�5�|��5���&�:ݬi�Zדoɬ�a��q	H���7R`�N�hѻE+W����R�i{N�to��wE`��vƟ���5ɢ�h�h���	*?�&�X;�I,l�E1��a���v`��:[�~ɻ������إ;�����w����XZ��ӽ%=7iݽѴ�\̹�S,CP��:�J��xȺOÆ��v�t�g��ӆ�����f�V��(�,`*Ȓ0���Y#�ix=���� ;_�ۧY�Vb��j�)j��Y�-75�I>v�L���p��x^8�P��خ�{y���N�����_mu���έ��w;�oy:/�]������>������0t޺9��ϓ��;/"��9x5�r|X�N�Z�4�_ni�7ƞ�ZƗ�>����e��YbfX�7��BH��-W�y��j����5m?f�E��H�BCNzΪ�,A,�I*� 5��Z0�+������'�.����o^�2{���9]��M7���������dg{x�J�)���%5�zh����qc7���Ȍ�TG�C��>�%n���Z��3ԗqV�ĵ,�u�-n�a0��H�9��Y�3������1��P=�v͂���؁�V�%�4���6&�~ɒ��-�`�Y^	k�$a�n�nb���p��/�� LO`���/i�=���e߾��?Rk}Eܹ����v�c��eKˤ��G�L%�*fa���9�{z���7t�[Z�W5�ػ�GХ�r���@2GI�+��@�(�$���`�;���[�=pݍ�Z[V}��5��R�6�	(Q�)�AN�� ��/�7}L�/��ƣ�s{����-��<^�MC#�{��K��}g�V���3i��Mu�E��9��A��"���qj��J+y�sm���co�6�cO�r��z�{��M�����7����0��O<��:y���t-OV��� yB^�	�	���[�$R�ў�s$�(U�9�.��{v��c{�>�v'Y����]���v�un��/[�z������5�<q��ٞ�}V:�&�����ڑM'8c��f�]�^���7���/n�nX5oܮ�MJhk"	��zo�@*J�����#S���O��-�Kg��J����Ew���G���{�%��%��|��R�&�J�<�$*%��h?o}��_jz+�}��=��?����	u���Fr:W\��r��������y������������4[�n3>1���~��4*��v�H�"YoKRjiʪk�f�Y,�r>fbR���V����v�������	m⼗��2Y'3Ꮄ5%^��P$�K��������w���ջS�]w#�����,�v��J�뜹uȖ��Ӌ(au��͏��Q���،iGgZRkZ��pn�����v��Om�ı�Gi��qy�1�  �h����W.:^����i�h�m�C��hҴ�y��"��Y��w� ��V}�W`��tg\kZ'Ye�l�!1����Ʊ��=��n��2Һ6'Q�X��-[_�56x&��&&q�J.<���F�7m�^���"2��(\; �s��~�.���.�}YY���
x\Y#�y���~b ��#�V�<0n3uG�}/��Q���u��=�����W�:����z7��ܪ`�N�#*더_+W�*��q��݋s��J�P��a��� ����}0P9��zU� ���yUB�9�=���#��� 愙ᓪd�f]j� �k�Z��W���ճ��E*T��5�bX��X�X����! ~�}����s��뗘�Y[�nо� ���� �����DSJ��C�fm���X�UQ� S�G��H㳻��� �c��Lq��U�I`?��� ��ׅ�����?b ��y�:K"�]Y�yX�W*:�LVf�#���]@�fF�]�r�wP�j<��ϛ*����� ���3{p0�k�-Y|�J*�@hW�2j�l=	�� ��޲Gb�s��G�~8� ���-*XHO��'����w�3dcא��
��H�g�I$� &�#s�=Z�f���y � �� oyw�U���Y��L�T��YP*���FS�>ͻ1�(�rI�z��yk�j Y}Nx�ϟ_��`���������W�ڿ�$Wۊ ��ۓ�c��?�UT﫿�N��������� L��� ,Fݮ��?�����=�/LjZ������8�����ԑIbyn.Tl>Am� ��]�;�I'��������� |�]E�p��?���}� ��=&.��ac,��l�L��g,�[.'�������veVNN�}Z�A���}DR�;��� ���ې~㜫�P[�m��<p={}��?���4���umC�W�ă�h��T��%c���#L$�K�i��L��p<jn�+fw�E�S�"�BȠ� n7Z0?��+�`W�����4b��S��Y�9��*�ߕa���3'�s�w�ް�:����.��{'��~��Ǥ���;r�HtWzr����S��Ӱ�����:b�R�6s1i=$���cMmSo#�:��oG_�5u��n���A�@�Gz��:5�hj7V����q�^lvK8����D��U���h�(=E�3�Y^��c�Ϻ_e=��{��=�����}4���{�ڧ�;+#�=-��F��y�.��W��-1c�����,��uh}7�Jf�N��uۚ]ʵ㒭��;V,�4���q��G����>d��
3�o����������F��[W��:M\�`y��i�U{��E]L���RPD���� ���?��rn�����Jw[����h~�zS��NW�:�#�a��Η~����G3�?#ː�i��ЁKh��EQ�v~1z��Vhu��5M�yU�K����t�0g<�6��a�VC�������`�|)m>�V~f�mr��[U�w�P� �B�VJ�1�e�.">ь�ʞ�hx�=[�.��(лuۮ��~/Icw��ڧb0z��?R�η�e�2�}��~~,���vec_��4,���W&���YS�zeҞ��� lu�p�rKV�慍"MVJ���L�Lz�����hԩ����q �#����I����:[�k>IL;[[�FP�i^R��CY���k�|������3��_���_p=��K��e���w�-s�u���ϵ=5�k=��:gI���{Y�-��^���Ȗ�<n��e�6�O&~���>�=���3��/��Q�v=���U��z�}�S�֮-�	�[�����%
�?)�S����n���.��vF����7�؟�z��N��kK1��y�ۮbe���R6o=x�(�B���ױ���i��W�?L����PuOvu>�e��\���w}]�Xմ��������ƝMlm<j��Q��q�p3Uԍ��qՈ�SMy�=V#V
1P��߁�(q�Ȝ�(!�IZ^�v�]�Q���=�G[Ө߳iL�d��ly���>l�
�!{�Hy�e�"�����?t?J?s�m�j��-��_�}5�c��S���rtN��:�Y�~��.�ѳp��M1#Y�P�6�\K��5�n�t�ll��.�i[���;ӵ�ǤY��ά/\�J�
���ȨL��g�)�ONJ�Uu;Yݟ[�}3�;�旡굡��{̓xS,mO:J��aW�̅��7��C���7|:��S����ﺲ-��!O�{g�Z���������zo?;
���~�ֵTT�Q�yXa`C����_�|3t�{k�+�E�ܽ����^[TiٳRxcjR��;8+$��`�n��}S��;n��#���;4#i�-�Q֚x��ұ3۝c�9�B���pN���N�v�������jݽ�z�U�^�����j��T�^����i}��xh/�i����'Qke`�+�i~;U��ďY5��[Q}Q�����-�E/��3/pd���#��c�ja�r�6v*�Az-�l��T�B�U4U�� �C��E� 9��h��W��x��[�/���wC�s�p;BzӢ���MG��Oh�������Ѻ��r�� �wSMm>X�1���5�)ߎ�,w�7���#J�՞�I�o�2��E�5zM����ꑼ��A='I�{�A3/�k�"��&z�Q�_Q)Wضlmۚ��]�J��L��I\?��Y#Q*װ�Ӑa�(]S5�������v��{�ԝ���^��:�WVuV�{pz���B��}m�j�v����`��bj8��qOr��\��=��;�[���6�}��Ea���D׌"X��j���x��$���GosD�(Q�]_[ݝI�g�������w�k�K$��7�%�%	[B��B����#�z��~� ~�=��?�v��ϲN��=��u�zO��kG�wK_�]G�e=�u����qƅ<�*�>V�q��N<�n�>NX�V�ok���f���xVj���D�4k3��|�FQ ��.|�!B3�.���[#Ou�KZ��!�Gb80�Zx���'5U����Bq�_�gu�#�}��oAvGI�5���������޺�]��Ӷ�u����n�ߡ�p���7H�q��3�o��^��v3�IյN�k:������s���b8g�f�@�/�Co�'�9{�q�VO֩;Ɗ��� ������!{��*^�Nw�f���<S���$\4�v�)$��I�9��?Q��7+�gqz��~��>����>��Ө�����ej�� ��C��gUӴ<}7*b֪� U���埏��D�'�K�_Z%]�wft�K��@5{�����2J��֊(%"U�|��C�U��r� �?�}Z�KvuSS�����=-*�b`����O$��{ة�	{G��K�y�/]��gW�/�}��.�њ���f�'NSY���u��� �-���+##�u̝Qӵ�C���hgO�8���:�N#tY��ѱ��q���-Ȕ0~x��7q#���SY��	q
�0���;���HP�r ��=��A�����_��#��3I�OC��z�Ӧi���5������Z�JO�*�ԇ�Q�jV"cM�w���j���!W�C��Y���{�R�yP��+`��=(�������������k�I��#������w���7E�]��w�n��;C�=�֭��]��5�s?�=���+���I��^�ێY�|}&�����z��l��*�"�
�y'�<��� �x�G<�p᜖p���A
>��?~>���  s���|�s4�3�~�z�/���������3''�}�ĶXǞn�91�l]>������T&4�>Y* �b������� ��<py��^� ^~<�������n������;=��^���������gMh]G=#���K�zrھ.��uMro��=Pu�͵o�3p�����Fvhh#�42H�^�D索�!ύ�� �efÎx6�5 &�(̪�����gF(�H�~ݼA�1� _�j�t�%�7K�Z�Nj}7���=g\�;I�Bh�X��/�Z~�E��c���1�%���Z�ۆ;�5h/S`�hC)`8U)
�x��M��<r���y[���#|�z�=�R=x��D��2�x����w��������v�[wc���u�qZ����t�K���8�=�t�NN7����=K�R��f��~,_ԍ�y�XPbx���Gs��c�=p�J�d�D#���< O�	 ��׏�'�sP5�SO֪�z��5]KT�^��j��e�G;T�ڙ�~��g�~],��(��ۖ'o�]OR[*�W�q�����^� �]��L���O�??������P�_#�ד"p���,�b�DZ�;Ou݁#��ے}fK�i��%��h��7cv�W�d~�����9�)'��	��\� ~\�=/���Ś�SW�L1�HdQ���� `O�6;�����Դz�'Q�ɶ�*���S������?�=g�=FmM�i� {��y����t�#����W 2���͢����m=���!7����Au�}]����O<^��8�?��dm��,����/=矷������c���Zajy�F���G�ٺ�Ů.����l̕3�� �;��7n��hۖ�z�m�ᓱ�y~�����~Ia�5��AV�5��9�~	�����R���q��wv�w3�!�/�4��Μγ��ci}KP#������X����96����_����\�V�̖ ����ȏ��8�kU��o�!�jD��T��N=�1ܾ��y��_��P�{�톉ߊW��>����z��im��k�=k�GV�K�.9k������7���N��SzǶbk_սO�"��04*���p_�n�?s���1���쭾�����:A�*��i3ʶX2�	H�!/��'�{��^�fi��.��54�.��[�k����ig�x�D�bo�����bx�Ly3��@��s1������oR��U���!�yYZH�Q+I�M܊�ԀsC�t����}o4ݽ��+�ܽ��K���W�aڴu�L��Y�LeH�3-�W-~��gi��/U�^x�N��K���y+��� M�W8�E+�	�HrZ5Z3�ƭ�nnf���Բ�л#��w1�+p�O yc�g{o���f�mKvmOH�fU�H�K<�>fIZ3�2�
?w(��oY�����\uGF_��W���5���n��ܞ��p��K�:�o�}G����E����<t���X��*E��h�V�ml������-�&�%�B
V�[Jq��Z栵`�J�ȋ�ic��|l��cz�I�nMϹ5�eT��Z�V�'�2G,�(In�1O*�J���!��X�oGV�b��J���=�u����>֝G��_�~��}���'UӴs���ot���>F��s�b���8i�����Սɧ�SD�=QС�tm�#��0V��.yc�E�$k�c�:R,j�{�״$���W"��WP~����:Q��j���3q�f���/I$ʚ}S���^V�:Śl�ıJ��8Jݿ�N`����s�I��1���F�zNM�yQt}g.k���־4%l��8�6�o^�V-Z�A��n���r���f9�i��>v�cb��A���~��k�GPd�����ښ���2�GS�$i$���R�ص�'�p��dv���pM�_,�ە&1��UP��!`*뷘�߈��:���F6X��@�FE[
�;�<�qx�5�G���Hf���<G�0B'? �9�'p�Q�8鼘I�h�:qM��!�}�X��!"y��'����K0� ��[�n^2�;�n�A�o&1f��&��S�L�W�fUz�@ ��|wؓ��6݌���S���2'4�R�]ӟ/��*-K���~���|D��Yiy�lg^em�Y��F� 2~H B�1ˆ�m%��7��Ew;�����ŋ
�$w-����J�lQ�u����g���&��,��X�/���D�z�ViD,q�X�nvDW̬ϷTFr� Ōc�ڭ:5�Fk�iB��<O�r�-����Lb�-Q�\X�]��[c��~��s�$�P���� vcT����2�ځ��V�� m��a=��\�@&�������D�� �W��d /���\��IE݂��f1
��b�iS�K�$��|��6A�ݟ�AR�>�c2-7u���l�Y�U����f�?n|xI}�}1��Z��Z]�U�S�����t��I��w	�����33�����R�-E&����J�(�;�~�@�`v,c���7h���Y�㌌�e�&�\=��X+}I��1%�݌& Fh�Y����|��Hx��h2�����3e*~B1��9d5�~~F��+��P�J;����y�Iʇd#��Y-[Ii F/ļw/uL~	2ۉc�`K3nG1W�Fe��w��<Z«T�9!DJG�=��6B���1����] �:o��oL��̙L��Ö�P�~X�H�ȧ�V�]ݓ�@ƊҐaI�X1�" n'm�v1�� (�ER�6QLb�B%��uI 
�������c*�����%������4��h��#�m����Hcf�#J�8��tYф�V3�FB�-wQ����zc�]�i�'�k.�K&,�M�E��ՙ������W��Ȍ�-��XυicZ�ھFD��8n�� wv;��1��yY��26��7�ifބ�H��!�\��119�m2���d"�y(��@~.vbW���4���@�lܘ�" �CB{H���n'����B��`.ʔ��<g�����Ugq�#�X�ggx�ϚN� $D��Wƪ���jTHlY��%w*C�f�f�Z/$ޙ�Q����R�.�Fo&۱=��s�Ƈ퓲�b򘌦�U����7�
[�-�c#�Cǈ�!ބ}��VE/AAz��x�*��%�1�	��@I~=�U���I���(HdT�U�.���-gŲ��&)󣆉��n��
�7�,~}6c$�x%�P���ru��N�� ��`� ,w^D)c)\4�h�!)VIxZ�`U"a�BLo>;�؎$��0�ˬ�4�8DD��ق�� c��  ����3�x!�<8�d�˖Է3B[���F�~��Ic+D����"�f�(wf(U�'��X~LבU�>���c�r��u�Z�l���?&L���	U@Ϳ�q`�9��-������ b�YJ7"�2� �l�*�v*��N�G4��Σ'����iM]h� W��� т�ۑ>��	���2"�
C�:*QkGF���dugY0$n���=1��P�G��*p�r��h��!��"K��0��iF�@�D���E1���s��,��B<�9���3��n1��s���ܲғ�XD���:BF�,_���D~\G$l��K&5(���6<A��c�Ef/�	��k���9�R��EzD�h�"c��̳�jfTدܱ���h� �&QVJ�D΄eK��'�6*�fv܂Ϧ2�Z�Ӝ����,εZc?�(I*���; Yw錎��#%x���~��2�YX�MU�oɝn ��T��Eر� >d�y����"���Ȟc%�E^�~�0�lx��l��
�
R�k�L��j���e�Iɑ�(� ���#���2z�Q�p��ڶ���v���Qg���ߎ�(��#d��2���M���i��Я�݇gT�K���i�*�b�Hw�<w*�����#���Ԯt��4��N�z{������}|�����u�������Ǽ���OP�tG4�����_��4���~�}�AS�Kǆ�
�_IP�O���J6f���j�Ώ䚮��c��J�R3b���h	��KQ;vHJ��^Px��u��9��ԃD�nj���v���
�A�m:���,g�*���^D<�h$
&����؇���m���>��>���e���iZg[u����\���MCGմ�I��|�W[֨�W˖66>.L���yפ�F�F�q$z<�_=�/y*�/)�f�p^4�k1�p�䏰�j��j���UKk�u��><O��)��eB�}K�����oݸ�� �n�{x�~����鼾��+�:�����I�<}Dɶv~����`�j�Wg��t�a85�{��S$�5�5�Sjͦ�F}S$�B����:?!;K^�C($� q�v��G�s|�i�h�!Y�3�^U#��_}��}�9e� �=�v�]��Y��]?^뎕�ν�{adC5�Nm��h�N��h9ֲ�fE���x�.�h����=�5������d��Z��>���${bib}PW�k �^Gp��'9��4�4�W�;�� �&�f5᚜0ךVR����m��Qw�D'�>޿KOq���?y��{�=��Ƥ�����ujt���2��Ұ����Y�,�����6��=0�^�.��X�X֪�I�aD�!�9lؒ(R=�Q�E����?����j�:֓R=7G���X��4�k�Z�x���:�}�g��]��?�o�߹�?������g�_@�B��X�O�S]��4>����0u�U�11� ����_�p�� ��yPE�R�{�_�%馕z��ݖ$K�j�T�Y��9dY��(p��!*�eN�$�6\�tޏu�sV�}�����Ң���F�+5�]1�Ҙ-D�����/���c�H�WS�� H;����w��Tbbu�����+��tj�X��u&?S��N�ɒj��|�Ξ[A�8̐��?���WpU�]r��u�����@�1r����O)�$�}`36of��%]=ֶܵ�5=JZƴʔd�th�iK�jX{Uo� 3b�ö�������ۻ>��/����;E�&��k:�Gq3�[��uL��+K��9��Ɩ��b�+�������=��[�H���������-�uo��
�t�fD�Z�,�'�ı�q�E³ʳ�h�}#�L���u�����H�Qi�KgR�� [o$R���y8�Ȁ�vF��~���R�n����sY�d{�v�J������} t�]�=Os��r����2畂���m]kN�jzXYd���"��Z[��Q���]=S�۶p��)o&��Ir"�٤�q��dO��<s��䙦1���ƻӻ��WR�u]{hV�ɭ��X�:��A<z�X���$"?$%l��g�l�[�CwϬ��w�]k���w�]5�|>�����꺰�[?�u�'^���j�T]�ǭ����U=�G�����֣�7���4�W2W�JJ�CV5��	T�9M�)�$���̳�[�m�z���ٷ��P��jةid6lN�^YS�0��M!���f����7��p}5�oy���� ^v���R����wC����uOs�f�9:?L�綺��J�`d�rUL�w�ϩ�g�dj�|�>V��TU-K<R�vc[d�e��1��-d��q�q���U�8�I���*jh{�G��V�R�#T1QY%�ʔ���7��P�2��O�}a��_���ˢ{׬{�>ڰ�1���j]!��^��s�������x�~���~�:ȭ�5(��h[#L�-�V=�ԭ/���}��6ޛ�mEVJu^���>EhE�>�y��bf�b�X�#2�Vw9�nn�^�l���n;�2������Y�h�$N---N%��hD��m��U�Y�y�^�z��?E�O��������K�uQ��@w#�5N�i�w�ZR��c�0I�.�\�ZZ�%"�7.r�M���/�S�з.�c�۲�����]̭.�9��>�<��� ���e�t�_�"-�u������X��BȎ��{:�SQ��|}~I��$x�Py����WT�Ư�v>�zkL�?y��[�z����o�ݺ��E���~���%���N���W/Sic<u��������&o��wHٛ�S�{�z���4-�V��F�ud�5+� �{�ka�"�Z�| *���ޙ��k����Ӵ�_^֯Y������3K��&��8��d�y$�y�>͈���u�ך/`����ݭtǸ���:jٴ��Dh��.�� �w�?Uv�r�2�N�U�����N�����ʑǓ.LM�n�KF�Z�����;8��b���TIN��<� �ȱ�c�-���Oj���{����R���39 �x%}��7~C������k�P����Ω�Ӻ��{�Z=�.��po�������m�Hix�����_R��+A��q|y|A�Z�ѐEjYd���	!��/��"�>��c�[�Y"�'Q�ξ&I8pʼ� O%�!J� ��0�	�O�^�z��M�MKQ�4�MC#/B��j���t��I
�����,�흖i�V�ph�D�Y�}������ '�8�Ï����A�UV1ءUG<��~y�� ��aC�P�z}�t����Nn�B�ڬN�lG�o��G�fR�O�Ӓ���r?㞍J�7=��� ��e���6� Y]Rx�m����_*�������(�������~?>���8�����<�����׿�a�SHz�F�E�y��޳!���#����� ���^%T���}>ǎ�H�!{���?o���? ��2.��C�� �z��8d� ����c����u��yx��������� o_1�E��%����}��~�� �:�ێ��5>�k:�6���}��\�L}#O��3?7J�i��B�eO�-*����� ��$Z�U.e,�}!Oa矺����$q���f�e@� ǻ�{K8��_��G�Ǳ�ulK3�q��t���y���FV?P�d!~A�m� ����VF����<�C�G��'�2� ��7���?��2����V8Tbg��5T����������#q��׶�(�y� ����9��M+����� ���bi�&\������4P�iϗ�'+bJ,Vk�6Ǘ~|�5b��� .�ϡ�~?��s���A�VR�?���?a�?|����뙹�>�|�$1�)Eǀ)��.x棈O��m���Չ�����(����I�>�� �Ϭ���������I�?��g�� �:�6�������AO��c�ʙ�fhY��N���+�	�h��f{r�����_W��~��jf~���KtRG1�}c���6ܨ�쵚r��$^J��sʖ�I}|:��m�x}�{�������oU�W`zۧ���=�͇Y�����5IQ�.��A�zP�YEM��dj�ΣPï㙏�=�;�^m[�Λ��bƅy�G�hej�H�؋����:J��8��N��v��ڶ��5�!�o$��ꎎU���Fđ��%��V��Vu����~�G���g�o9=��\�nH��b}���S�F�ގ������zӨu�Ա1z:���5c�b`b G]B�%Ǐ���/�tyn��t��j�i�1���SQ��U�,�����L�i�h+�s��wJ:3'\t'yn����,�I~],Dg��m�K,�X�)*t�bf��@X��We{��n��ϭ�[��{����{O���/�>��۾��� �iyZ��ߡ�깚Z�aj�S��ޡ�t��(�4�	�n��O��:� ����)P�:�^��=7O��k�P��p�2H�Y��FX���Nb�#���}u'��:%�>�ښ�\��S��웗�`���4�&�)gL����zc2A-`�w�I��aڏ���Ω�}�v���^��_X�﮿�S�:��pu��g+��-�n�Բ:{Z���OZ���ig�O!r����7��tM��j�� J���pn��5�`�f�(��J��:t���yYԡ��O�=����um�_D�Z�r-x/i�y�R撍��~��I�d*�/}���Ot��>�:#��x;+�=����fh}1�à�����?Pj�m�1��_w��yew�W�w�>m'Ӛ`�v���x���[����;o��;fQ��>�u��dBkEnX�j�㞾�H|ҬOjW�3O$�U�z'��?zmͬ:.���4�T�;w�{�B3�4�엄����ҩ�?pV}U��E{3����7�?j���Oe���]���zz��{��k��׺�#X�Kt�P�&V����f`��L�J�saf��;��⿩�rh[C{H�B�;��:]��:ma��2D���Kl��^�_TJǅn`�;gi���lŵ7>�RΡR�	��� �
Ӣڎi����>!�E1Rx�}]�����U�J��vzw�Y��� N~��e{E��!�XԧZ�t`��m�P�� �lw����||7Sդ�+��kL�F��G�$�G����}�N��p8� ��ϭ��������#g��B���I�O�@A?iٳ��������WN��z����@=��w�����]o�5պ�H������3��E�6eP�]G''���6{�i곶��i��|�rW��У>���RV��Zqj5�7��<�MX	r��h����Vi��_�=Z�lom���o=Y��$ڏm����5��v��a�+i���۰�����{��}��G�>�Oe���=ܽ/�r{}�w���������,bSU�𳰴�z�`R�ՠ�v���<+|>���:������z�j:�jo\ڱrQ�uI����#3J�\\)�,��.|AtK���#Ԣ�KO�g��V��jF���=Q���|a�9���p���������'��=��{�����Z{v��:�L���#���x�t���&��fa�� ����R}u
~�t�J�^���ޛ��rd���:*y-oL�O�>��"x?/u�S��/T/i�����R�*q�;�{Ǿ<��ӆ�X�H��iߐ:5���:��� O�����O���/�Y�?��wH�[wO��[j��MCN辬���JZ4�̸�-��>�k�r����@~:�� R���SJ�Zs�Ƃ
�Bi'�5S]�ͱ.ֶ��QTƋ/�+,������5�:{�������"��OpjmH�a%QN��l	�R�|�F%e1�v��/b���K��ܽ��G�m�Ӥ��ݴ��];}���=3�}g�=P��:N�ҙ�W^��7�q�#*����g���:ﮨn-ǢGCK�]�j��in�\ [�Zn,q���b?
�cu�6�i��I���n��=kY6̒׶��H�E<6Tp�yI����+������=��Gv�N��~���:n��%~�����az�
ІvNU5��E�I;���*g��&�i����6��:[�9ι���Y���J/���1F�� �Б�Y�A,`�#�}��}��k}E����mH��0�r=4r%�֓��,�F�+�0�z���{3���������]����{�׺j�?��PͶ����]Vg+�:~�U�=2��e�/��L�sתP��Mƺ��������*\R���/<�*���d��Fc�"(�}2鞗�m�-7� �kZ��ojRG����ܗhk/�=��3I'%��۟�k���q��T����3��K����W�p��U�[���Wd����d�%e��V���J<$aR
���K
��Enұ�+("9|�n�~�J?�3(���ڦ��rr�J�//� �>�1�W� Q��~��O�k�1�s����ε�}�A��N���B�I�߬5�W����5<�]AƲbSmE�<�����+�e��J�V���9<��8b�?v��1B��y�9�W�sIӖ_@��Q� ���YO��^>�ס�G�w��笠��ތ�\��N�?������w�8Z>kt�L"F=9��y�P�5+��x��ԵF��ܖ�K� �?��rs���<����<� p� �Η����g��C�����f���wE�٧V�?k�l�=�Ҕ��߸�w%��(ϧc�B�����4m _��#UI۴	f>�����
��ny�ɷ_�^�-%x��U��`8Q�$���n��8�Y����w�eӺ�����r�/��:����Қ�6E4�
�f��U�Kf�x�gC�*���g����@�* �[2N��Z!�����9v�or���}e$Z�iY���G���T�y(I�Gh'9i��f]���X]��_�>����e�e_N���g���-gL����辀Pe��Jr[�;�u<x阊L��f���i����U�$��R;�Yx�����_���߄���i�
��Ā��\�!�NC�}}<���������w�����螗4�OgS���-_?�5���T�wP�O+��GH�yo�\�`i�s�]GS�bW�?q�#��������R�h�v���� G��9��o�͇�B�w4q�%~A$�!x�Q�� =TP�Ӆ�0��� w����ϋQ��T�_��_��F�Z�:���:���P�� � +@Կ�G��� �� ��4��23�>�� �O��� �PNb����q�����?�<|��%�2�����@�?/��g�>>ޭ�=J���)�p�<�$������ �WשZ�2Υٸ�@z���������F���5u�v�GfP�]�mE �A� �oj:ջ��SQD��)q�p���������N���W�G �o~����� <��鎤���jZ���8��2f[��e��~����� o�WK{I29��p�n�b9����?ǌ�Ǯݏ��u'�I G�O��� �k�[�~����:g7Z���k����y�Z}a�6|Ժ�1����<C���V�*�c׵MOH���κEr�F�cVg��cg��}���fI�R�z����N�`�U��T(���=� >�z��3w�@�ҡۼ΀�}k�:W��kZ:~��t֩���Y��u�[!�~��^:j+ddD���R���p��Mm;L֛Y��ؖ�ȡ��1/{Xy"@#� %��U��Qo6����jZ���c�c�d��Fp� �Ǟ��	�(���3�W�GE{X�1�C�4��h4�܎�aa�?�-O��:�C�gj������G��.��z���$2qu����ځ����G/�v]7�hl}Zm@;OP���Ӈ�����p_�i�YZ��k3i��	D��]e�����s��4�yn8'ҷ*�zQ�n)���*3��c�N�4��1�:V�y�����i�#.y�;K�#����ޚ��i��?�o�mD��.��zl_��=Q�e��t�"���N��x��)6��%Fw�v��MG� �aC��m�.���}2�?N���IB˒9kQM0fY� 9m�Ss׫��N���+3��`Ԛ�t�����r�#���x�i[�'��Q��A>�wS���M鮪��z����F�n��u��<��u�Ofw�D�5Ρ�ֽ���hi�X����|l���ȵ.�l=�����5������5]NPkSӔ�j� �uR��J�,2	�:!�5�����]�j3��A;R�y���:�It���$?7V�*��T�#_�,�wrRF�����N���;��>ͽ���[�é��Q�uop=��ι�}����`�h���b���N���MJ�i����?[���q-	�ڶ4��:f�����ֺ��*Z6��aI�Яj�Y���!2I�5�Ֆ�ф2i6,�I%�Uc*�����i��'�]?���NC ר�SU�V��!�kK�Z<�+K�!բ����	|������{�m���7G{h��.����Ӻ��׺�F�Ĵ̾���XdϦC���ն�Ji�4�I���=b�z�{ӥ���ۏR�Ҟ�K�X���uuY��-��;r'�D�*2�ݤ���'���lΣ�:6��]�m~N՟,q�)�S4<u��5e�:��>B<�ø��	���꿪wz;o��V�ѽC���������]s�Y�i�J�?�b�Bz���*�X�y呉�k�@�k��Ď��5D�ܲ�%I!�x�� `�ffI�V](�yW�i\������?�gS�v�˱42V���eFx��,u��I<�ܒR�%�4�q�� ���_n^����� kߩ����w��[�z=:7S�0�,�O�5XkT�sc~����>F&�ؕF9t�^�Ԏ8U�� �-�й�KU�擲�Ԏq~�k4��#�cGJ)�	�Le(��*g-���z�Wi� �ձu=��t�R�}K�$4r�3@/����#�d1�Ѫ�]���׺WW�IuoKk]!���91�n~�ԘP�j�]p�R��j�X�M\jUJ;(O5}P�|R��[��,jȶ)Y+��YO��	��s��8�7;J��jò!%;�ƒKN�xn@��3@K���X�H�V�e|��}�e�w|uP�:�2�)�^T%+���,�x���k�ݼq�C(�h��T"�"�����
93�@��1`��Oї%T��X����9��X}yp*X��s��<��r#QjPq�33��g?���>�NNď��u"aU��� ]n'g�E�ꫳ�1�c�vc#�Q���a�=��7�V��JV���m�<�v���1�cFV��gX���K�6�t�"�ʩ�fP�Gث0~FL�Y
A&Fm�79�Ep����QEp������,c@�XAVՙy9�p�t>@FCll^�S��O"��>C9���&�Δ���Fq%�I�ɀ5�4�hW�R�Y�>FG0<��֋<��q��ޙ!w1�� �Q��Pn�������]�i�|�We��s;"l���7 )�0���p���*I�kuCJG�%��h	R�Q�3JD�u��L4�L��# B��R�Vg�y��r`TP�6^ZXeJi���<G��W!�2�(��]����b���ߐ�A�NP�A�+����`|�@��n�X����T�7�1�t����Y[�x���W������1��,�)?8��|W�0Wv�1&��I�,Ǘ�1cf���^��WĵN4���'B UV�^�(��rp<a��Id6d޾><z��(n
_�M9�;3.�	r�@��l�!�ȧ �$���mPI���	�(���ޘȖ�W/̯F�IrJ,͛�'(SnT�0��&μ
�c$�Q);�e�c�$ǚ��[�SVtTߑ`5��`�e=n�E�H���Q�Ԓ
�:|��-��r}1������+��J�Ƴ2�ub̨�ŭ>_'ᘐ���Gǔ�'%�R�>�LM�F'��&FG��g�r�B��'�M�Q�i��h��35�����/&�����;���I� "�#�gc�;�W�E��:>����1��R!UM]�Z4�޾5�F�Tx�?���#�%@c	�h��?pڗ\J��39��VI�`��}�*��oLc[��θ�E�Iӑ`
X֔�6�rK���~}�*ª��%&r�<@䅋Q�EqAe�O�(�Hb�����g�R��k2� ��\�Rh��8Λ$o�����w�������C����n[��^Gv0Y�!f� ����4p!A%�V�%4ݘl�����2��y�[Aw����e�E��)�݉�|c�-�Ǥ����|�s~qi͊@y�C4J"�㺪с`L)$VZ"(o����Pm*2Q�U�
�2��o�%�:�!�_�e~3	U��q4eO
J�D�怍�	R>�ī�3��R����<�U�̲<*��Kɶ�[��e.X�	H 8b����o����<����� >��aIJ�i!��>`�^����β��m���;bŹ�@�VQ�ǲW�`��K�mW���"�$��aP��f݌;arg.,���3`�Ɍ�Ȑ~)o�}�؀�(!��
�i1i
:��G�s�ԏ*�uV��v5~A�|��1���s��h|�9�:��(	�2şr�@�P�P� oŌ�W;�X�a;�1w�G���lfR��B�����X(��^&Ş:Ҋ�'Y�@��)�G,I-,~�'f2俖Rȳ�6�xc�Y?2μ j�nw��P��q�����2�q�EFj	�I��K��W�nЧ.3SC�}�c�.ag
����"�!�:��a�G���8������*� ��)QH�[�4Q!)�eY�H �ݶ�c���G�e�= �@�g����а䠕GD���=�7�0�F����;�糥���/̺�C@�(�C�Ld
8qD���46(�����Ҩ���"$\��0ݘ�Xə�3j���4SYj�I�U_�_۹m��q(�ܳqȯ����"M��Z~:K�j��o��oɷ7C�#I���5�#0%1g��������ԋ�UV�aE�f�ww;\4�Q��4�sa�T/��{\�=��8����im���{g�'X��'o)�>�� }ps`u��2j�w}=�u�Qv{��m�t���%��������<% �>|�β�Zn�����q��K������\=C鵕�IcI��n�卾�*��,�DG���4�y|:��V��,Ԥ�U�9�o�V�k��2'ZY��P5y�o<2����{��
C�������B	��:�HjX���UV���z[����L+�1�#���#=Kp�|<u
�z���/æ���-C4q�{
R�y����;�8�x��?���ܱ���������cynRx更�$ұ^����x�
y�{�������>�z��������<�!-�=:�?�.s?37�����t�(�����Ü��5C2�}� �l�w����u��4�,���'2��#�^8�y�/���H�t��Z��m��i����X���r���M4��A�<�hU=r�φտD�zz�k�s�N�urp��=K�P��j����U}[#/L�� V�>7��U�1c��ɧ��њ�ƕKOԠ�)v�抜 �֎��(J!p#���I�]�	龷�j�d���Ҕ���yٹ,ZܕL-#1������2q�9� ��}����k�����>��7�K��W�N�g��C�G�:k'R��������L�p��p)�Za�+%O�����]rݚoT�G���;wV�������v�����5V�*��h�c$׳:�������?�o��m�4-϶���,/�G�|-i���NʓB�Ibx|I�=y�Xe�M���w��S�j��zgq��Ծ�,k�]����^��n���=OֳzsG�d�ӚG��:x�^*������M$��|4X�f������Ӵ}�nK�U��nޥf#P���!�2@�K#�G�%����?�|DOk�}0�Ʊ�n��I�<OZ�-9d�؞g�,���|M+B���W��ø?��.��ctf���ڦgwr�s�|�C'R��z�Od�Mi��Ֆ����':�G�nz��H.��uGL�R�07q_�E�2F̲:UUdskw��B�{���P� {Ҷ�چ���j��:U��N��3��,�6�̆�8�I g����i���d�j��������=5���{u״,��:_RҰ0�N��33��4�����*���.��F��Y�R�?K���W�&��^����2=�$��|��C�")��2���ʢF��Ŏ��O��H������EV8,�U�T�W}:^j�+$4i2J�d<X��įe���]����g~����~��{�jK�.�{��<����|9��ޭ����KNM28xs�81[�6&�d��,���&����GR7 աڶR�:T���fR���:W�*"H�5�%��v�P�(5���Z�Ov�i\�Uf�b�БAGL^ц�rN�J;F�K+?2��l)�k���{v�]���Y����׳eӝyخ�v��M�g�z�Q�A��gd>>��6�'�����b�d�-Ά"&�?��z�Hkm�>��N`�5
w�V�"u�V�R�;�l&9�$��ݒ���6ޝ,�$���5[:]��ޥ<4����P4�gF���+(�y"���`�ͱ�go=�u�Nc{�d�k�]]٨� ��W�;�n��|m[�I������Q%���c�l�j���1�?*8خ�����n�ӣ��n�ҍ��Ϲ(E!�F��m5�U�~av��ة`��H�rِlΪ��mQ�u�d���S�I��$X��u�i��4���WI��*�
M\�9~W�����?�~�Ի��xt������ɗ������s���U�>&��q��;���ղ�Q��|(��4�yf�%'�c:����y���/A�6��t��l�7�
�ı�r�VXU���p�c���)P���w�;� Z��������gAR�D��S���ec�H�ee��id O��=��� �k�����i�����WV�un�ҝI�:X���������е���ѳ��_O�z�φnM��z�dUf�"7վ6�����7�ѧ��9�iR����r;�M�I$�KX�������%���v}�h]���&����Q����*�E�;ҽ�1NB��3�_��4���{�Ҹ9���������.���7�}?A˖��]9{�_@eW�z_V���
�GZ��tځ�x����X�f�z��$��k�Ѭ]�\�]5�X�)�p�?/j?��E[*��2��y�W*��줢���U�aj�A2�{�go�R~Z�ى�u�x&2
G��� �=���~�e�� c���:KV�05�3_�zwS���K��M��t�6�=_�2'�~;b
+�+V�%�ԯ�wB�N9�j�J���Iӑ�;_��%Mt��fz�v�֑y;}�r8-�C�yR=������P�Zj��S����W��3��L������Z;��#"�o�E�~@�j�(h�Ɛ�G��@�v���?'��<�T�^ߑ̫b[���O㏰�}�n3��W)�^��GT�^d(P�� �v�������G++ڬA��������$hO,����.�4�R��kl��-Q3!Ld��5 � ��;r�؂�����~^�*�D�������=�G�?���z�=�p{���~�A���?�����05,���cL\�$��R��~%�� �oT�c�iI�#'��e�}z?c��e[Bm)�[����?9�szS4O'(j´��9�x�W�����)S�Hq���R���5���p�Ͽ��s��1(=�erx>���ǿ~�^����.1Җ(��fJ*����5�q�� '� 'ו�n�%��������dr����sZ�͸Fv_��c��m��� �����:����z� ��}3���gh=�dyz�T��SM�s�.�����'�i�������^�Ze�]>���vZ���4M���m6����DI��)�cer�ұ��-����a�j�G���8O����ޡ��.�S�����#���a©���Bhڦ�L�m<|��dIq[�Z��!�UvŞ�G�"����X�bx+�}� s���y��|�W�@����Ͼ?��eu<�Bc�(�34_!�P�"�Ȑ���o���-�\�Zv�
�S�?�����s�����#zo�� L���v~���|\A�[hz�����lC	s�����&5�bo>@ͷ����n;P�.ռݍ���+�enO�����ご�t�%y,V��,����@nH*~��>���~�{���;���n��}"��n���4��w'�t�uo\�J��7oz�V�\wZL?6T���麮\SǄr�B�7M�;�e�q��6���b�;�Q�g��'�+��تS�� ;����i�)нv��qJ�|��r���Riy�=��@�1P{Y�{����9��t�qzo�:� ��3�9x�2���8u�kp�=0��w�R�,mO�4��>D�q��k�erl�[������=��m���B6յM�T���E��n��ZEQ`IF%��f�ꮥ��a�i�,�������4ޟ�4h]�,w=i��H���lؽlD�;���a���l���*Z
���+7޷�������{����:��ݼ�u���Mi�ػ�׽��>tzc��s>�vu=c�2GQk=A�dGTl ��R��k��MZ�2i�썯�h�~T�K+�Ki#��(j�l١���d�����AC��+� �R=R}׭�ڵ1,��t�eV�>�6*���4b8�j[:G�׸g�އ�\���������	�-KI~��˲}��ι�ol��ҵ���k��擫���Ժ��MbY�6����NE*ͦg�1��ɬt��~��7^wd:��$��?S��u�6�f��;/<KKs�E�x-G]]�2	�k����>��G��ޗ�:�J�ݕ��bM�6K�%H%���Ȓy������jyT�����gg4���ϰ���ŭ�YԳ����o�'�>�e�V���9�}��uMB�^뻳�M-F�Tz_T���IZ�G!��:9��wfn>�l����{I�$�����k���%��f�EG�З���q�k�_��f((� �SV���v��45�Z�X����Ɠ���r٘Zy%��H ":j� ,� Y���:���_雯{��n����G~;��]��{�w�������.��hVM:�=���mG�4�����t<,]2�||�0�I�5�h�d�A5���lhb�'�PҴƭ���l�o�,�D�<�c�nx?B즷�}��%�wL5�k�����.jL@�?4q)�,u"	fe���O�~����#�=O��`����]��� G�}�ӻE�.����z����Һ����?Ǥ��4��?q�.I?�Ž�nzC��ӏ��[s�`T�wm�/�Kz����!�&�H�Lf9��f��W��juX�?[�Q�v�6޽X]e�&��4�WuI$_�KV�2Kdo3���y؎����G}�v+��~���v�۟[�%�yٞ��>�t�-N��u�����ӓY�3�'jeS+�� ��OY���.��3�� uo���h[thuG�Ma������X���E
�e��m$hU��,sҺ��� ����;�w�:�q!���xb���cǘ��
����ĬB���M�?k��5�l]�?t_Rt�Mu�_n4�uIu�������A����y��Mv�����,��i[���6>4���n{�{^��N�SSzցY�N�O�Gl��+�|o�Į�u�@�D�-M��ݭSJE�Z9L�!V�h��+5���'���I*H����}�wG�;��������]�������]Y���wPe�F�2�>/s{k�5������r�0��a]c�g���t2�ι�N]���ݿ�[k^�_��k1� �D�v��Mp�*y)�^>�� i3�]x��Ewf�.��6�;���it��3^Ǌ+F�5�E0,#�C�;">"�5��w��'�N�v��g�mk����߹�^Qh}E����^���s��?K�ӓ����JX8gZ���14���2vwMv.��:_�a�z��i�IRB�5Gr$��dy��CyCTw��;[�S!�#x�.�om��u'yͫ��S�#I�YjQ��<P�H�֖P���Eu޿HW·{��%�;�߸]G���_�r���X})۾��=�k���[��t�c��y�}�yi���F���Ƕ�ZzE��y���-��N�����}F���|̢6�%�,ۍe�h,F�5'�bS!�N#������W�Zd��ht��񙢬�j�I�� �9H�. ,�ƍ����sz[�x��v�\�/u��z�w:?��qN��Wj5܆ө�h�;�8X�lܽ^?��L\�'54�����������7X�>�ܰ��WT���P|�j�-ʓ;��n)�^;����$s��Q�G�r��旲7�֟fʴ7����tͧ�5b�!Jr��Q$�	c�)�$�f�H�[�}aL��>��������r�:�D��p��W�n��#K�����nr�>=?�ג�P)���� :�6=����}n��L�j�[��_N���$�e���SN���Cq���QEګ��׹Dm��������{����>Ҫ�b7f�nZU!�$��c��f�{��'> 9���o�-�����պ���+��}���n�L�L�5�_����Դ�KG}5:nZ���Zf�W\iy�9��Ny��z̚��<�%�,H�O7t��c+����r�~G�n�OQ���&��T�(��E*"o$q/b'r���)����]��_B{������c���h=/��uv���f��o��u=C����:��Q�W�Ie�)\7�f�<T:��	I`���Ve�BH�U1��?R��k6#dh�@f��(ݾ��#�� �r�?@�� �� �O��i�S���Q��t����Mo��w�:���i�����DԴ��������P~��0SU̔��X�J5�9��	��� �㴱?v*=r}{�y#��\x��
ģ�I s�1����}z���o~̻�����w���{W�3�_/�}�w8�M�u���D9�]����>���C7�oś��Y�S�~b�{R�R��.��rI����L�=��Q��@�Ϡ �~��������Y�'d����.�uWItOLuWJ����ɓ��W�=���-c.M�����6���� G�Ȗ.i,hm��T[v3^���,X2!f���T~�ￖVbHP����Yg��G�[��^Cs��Hp>����0?��?��=����_L�k��{����us�� �Ӵ��֩��d��.&��h�*��1�f\~9�m\Ghg3�SՏS�^�l�$Vy[��g��	�%����Ӵe�.D�]B�#�v�~�6�]}����9���Ժ'�$�zX�.����)׆m�~޽��D��ЫMa���ƙ|��"}9�淆�ԩ'���[�%�����>���q�v�����c��#?b�h,�,J q��G��_�H ��?;��^��Reu�p��X�.�֚��Qk�/��e�I%8��`H�6$XرU�4� �?�!��� �p=�������'
���������<m^�]$��T��]�M�qr�O�������i�j	�fG_�������ymk�To�e`>� ���~�3O�L�dAQh[��㒇1_�;�?���͚���g��:p>� ����f��7^?�_��ߞ��wGѠ��9�b�"�!_{R�P~I���Y�Y�A*��w?���~��??|�4t��.��p���� ����S��\=%l; ��P�Kr�����|��bI!�'s~�Mb��]�"�3)�7�s����i�I�HV���� Ǽ�Z�~�8Tˎ�����`��o��VvI6[�+JlA�7�����+i��n�s#�O$� �����Է��$�������� �,�Y�(����KU���ŎV\�(�q��gƬԡ
C�`?����ic3��(�nJ�N�� ��S�̞M"���k%�q�q���~�f�����>��ޒ训ճ��j�?��tP���C�io]3PԴ�_�:�&w��ΚV��>oWi��ML��n���z,��݇��o�[qS�b�x�j��m�)���$Vʷ�:Z�+-ei8�*�;�O����h�.�RJ�I��W��!�#�Bw)�嗙�¬Gi}��GD�?��޻�ӾｵG�5Z�����=;��{ھ���zGNw/�;u�iV͇tz?F�u('Tv�'P�D3�5�i0�8�"}�te�.�Y�ɵ�-
2���kybе�˧���I��i�dW�9�D&ٍ�F����t�
��5��X�=_K�X���fD&�����v����O�#�MY�`{��Oէ����Ε�3=��N��W-����tn����~�Ҳz{��kQ�Mi5-?-z��*d�+a��+U�3/Jc����$���n:���%o+j5mZ��0�'�T�E�(�N�=�4.�ŷ4���^�x� �VqU+ �'��71q��	�y	�Gn{�ߧ�v;�ؾ����ۗ[��K�Z�s�΋�^��])֘��NV�~��zk$f�/vV]zXZ~����q�	��ju�ϭ���ػ�A��g�_&����Yʒ-����|Pik�L�9hcc �Xw����U����5m�j=����50�d�h����gR���}���2:��4��/{�W�;��i���Z�d;#�=�wKܯ{�Q��=���v��-G+���X��%Ƌ�N�[��^�{Z��%�3��W���Π�7��q�����Pɥ薤��>͉�Z�؄�}�uEu׮�j�\��N�{{;bب�w�Bu�5�qX�l	�0������nX���z���;�1�U��� ���n��7��GA�Ln�����q�w7�Ψ��j(��0�cs��P\���֝��ԭ'�/ouQ��ЭӤ�
�_,n��2.�,��9�� �ZXB�n;���>��xֶ-�[����J�y��2H�k���8
���2�2�xho��������ڽ����G�l�~��v+E�Q���XS�ѳO�Qs5l}Q�b�$q&կ�&1^�|� ]6>�ܻ���c�:�5
o��N�����N�^.�v@#�a��� 9�?�5���u�͹�-6mǼkع�t���C�����ƀ��$I#3׏��W�s�F�q�װ�S�=��W���vߢ�äz������q��g@��5[=�����0���y��8 ߻�K��S���[�O�6���^�[_�jڭQ��	[3�$QI�"IY$`�"frG���5F>��[f�ҷ^��{����Z�r�Q�v��4r��E$��謅�P��3���:���};�>����k��}�h�9��]�=�N�j���p!�u�GP�%����j�1f�b[�hJ��i��_Y~>)t���J���_�B�M�D!4��
�D�wM��1V�˝����GÆ�����V.I���#�i�Y�	�4R�h��M��+�s~��i��#I��폰Iou~�;kj]oݎ�NZ�"cKD\O�\��[�'.�LT\	�%�# �ts�o���w��n���Ӷ>�B�9��"1�F�K޷���&� �E"F�dwv�T���.���F��{��˨o�/R�~�i�ƕE�1=ioG*�V$1<�ҵh�I�Pq��߷Lt�u.���Bx|�o������V�/]W�4e�JK�i�%��@@��K�}��{z��zE�d��3W�r��I�h�s�"t��H��/�e��3��]�E]>�.�l�f�A���U&�����M�@�B=��w�	�|�� `�&� ���t�dA�O��W�ǳ���b"6֍ֲ�~��p��d�cQ�u"��v�J]:�w�2�P�2����Rr��23LZ~�CU��2�w�LX,�8t,�Uו>��6�H�uV`�&RW����� ��Lx�:��6b�fC�@]�CE��~�[��p�|��p-t}[����.���Yd�gJ�!��q��e^���";>��'t���g�]�7�4����|��7Nj�:�N&5��J϶}^Y�.���<��X�/Y �%V��X�+($}ǰ=�����#��G������g��RFe�v���)I��[B�#�Z �|E�����o,��4���lW�,����&^ILf��V���P$��v��%J;2�9*�[Y:�Ɣf���܊����b��î5�EEm_ū񝤠���&��wy:�ؓ.A���1���R╳-����T�� Vm�*�F9b_�s(��*��:+�S��"'Oݛy����QKn��1�xe�x̏_���U�?�#�v7��KS���eV2���j,r��#j3�ȔU���{��O I���P��D��U��pfQ�*|x�Gf�Z6ʇ�*1
���Hi�-o��VQ�΋�iSY�Qa9�n�Y�R�o���蔟��d�B��⿷M��mO�^`X�Kv��nf(���|SeE�:�h�||T��,�ܾ�����c�[�0U������D**a�C�<~x�R6��
����-7<������W)�Y7���F� )z(Ve����<����I�)�! b��.�f ��e1�!4��o�x��0�M��d+�܀��e<�Ϋ;|$�l�%��Z�!U�[c�UM���µ��.�_��y_�%C?��m���).�~������L��X�gbT�TzQjX��$��|�u,bO�Da��m��f�l�{��$(�a5y1�C�d���ո��6jc���#�ǯf�ÓP� ���%�I�W[��V~P��F��6=��Y# G��2�Qɝ��c5v����f�Ǜ�4
�1���v��_��qc)��j掦h��Em�?�f�Z���wbF�w 2C�%]RZM�Ԛ�Svv(ª�P�n���J����)k�5h�9�G*���H�*1Y>�ӏ�l�f
X���H3����M~�v��I*�S΁��	_LcR5g��MMrq٨��*�H��� ��tR劰����h�K.D���drT��9����i �����?�X�߉�x�p�f��+�l7�/
�;/*�l�#�gc���doԢ$��X8V�v�ٕ��ߏ�1�qG��/њr�>V*;�%�M6
I��$�6X�fVj�Ҋ�o6�P��W�wU�n�F�ą�1�&w��zqm����!'�r~/�]�� 1�ƏA��LO�+e��Eh�ve#�,�ț����9��2�\iQxB�b���I?�'���b�!�M!�G����
�B��[t��ZA]w��0F� �����SD>wY�ADs �7*��`\�U�vL߆4i<����#�yJ��|\wJ��r�pW�f��#��� c�/˕,����5B%P��˹W���*�^:T�J�!Aje�����wU�؞_b %�$T��'.Y_�b�:�ev���g!���M���u
��I�� h���JZ���x�v��Q�h� .�1�O�g!���E
�7�V@&:��pv?N*���"�QD�`e�&Kt�P��9oޕm��?]��eoE�Q�S+�tz�m�,��U��T�*ʦ����1��G�֤E'�'�YU�*��y<�N\�8�����^���y�̓&U�J���%���7)���Q>%���s�k�J^`���D�*ƃz6�y|D9$�.>�ì��x����t���*Y��ܕ�g.���
U��f�
ƃ��
�s������4��,�T��ķ؂�2S��2���iBA&�pύ*K�ۀ�R[�>���}M��`�d���"T$�Ur�MU�A�qw�Q�B��r*3�	���;���8g�pt�o�� -�1�2 3t�o�-�Kxf����v����:N����LmKo�n�$�v����Ug�dGP<�deY{C$��;�:޻G[�&�^����{��~2�ɧjYk߉>�dbM{��4�2M�W4~�v���BO+�_^�keet���v�3'Z�N�gK�s�����f����^��k�k�'\�Y��گ$,�H�|V�8��8���e�aǍ�xlѮ�Gcv�m��hSm}�_�%q)V�9P�����ʤ�I���D�F܌�_ӋT��~��'�z����Q�^�tzK\��^�·Q�=C��M1�~���L�2�����Z0�L|����'�i�|��=�Gt&��)4�NI�Z�X{&�Ul?1ֹ�ONIG�̥�?r��7m��ѽ�o|��ͼ�ȥ%k�OAf�1-��V�Rd� z�u�?�A$K!N��ݹ�ӻۗ|�����zú7�{Cꎚ��o�i��s:�\���gR}���n�s���xf�W�O���f#�=!�����(�J�i ��g��hG�1�eJ�W�qi���9�Ζ��E:�mi�ua���ֵ�$���v֯-*�B�#I��;z�-���!�G��T{�����V��x�,���wg��1��W�t�'N�ǧ���vU�\	�V�xy�F��t��^z_�ŵt��Izm�v� �oIY��Un�#ٷ�fT`y|q��$Nf*��s��F:��G��.�T�����u�O�t���(Au�X1VF�Ψ$,�����;_;7�n�~��~�����}�{[�WL�v��z㲝G�Y:F��:�&F����L�fKM��E�0��%2�r��zt��;f��l�l��2��	d�Cl|���Xl�sަ��h�lBB؅$X�sޏL���F揩ƴ;�oЌ���^��p؞��,�ZN��x�2���^s�$����<�K�#��#����։���S�=��+AѺ����u��.�KuE<t����͟+,QqA������`FQ����K>�%MЖ���5x��_'��$�;[�j������%{3^��b4l��B�x����R5���dwU���힃�^�5wZ����{���~��g�c�~���4=K�z�?�t�6X�8�z���Q���;�Xf~U��#h������K��]7��\��u�6{	jݻ'���yn�1G���Hꎱ���	�߸�t�� A��֧�f���Q�\УV$�<zlI�ZI�J����
�+9/;3�E}����v[�<�S��O���{��WK.OD�D����}v]5�[KMOM�#,̶�rc�] �$2�������6�u�b|X�ҭۦW����K�h�[������ܱ2�b3�пrʌ�S�~��{�_��Ci�Rk��f�t�F��<�e��'h���YQE)x�&�ftI#:���J^��V}�#��z%�-72�G�t.�ާ�����D�f����eֺև���u�F;i�c�`���}���%N�s�ג6�)��I5H8�!xR�-�;Y�/�_T��kރ%�B��/W�
H�3'c�qIa��T��0gb�͋�7h�K�:GN~�ߩ��w�r�vV�݆�b�;j}a>�ѐ�t�ҵ�Ҍt�.Y� i���ΆFL�2ޣ|Olo�
�ѽ�N-F�9--�z�IbK�w���vw��8�y!O������>��8n�{�uOvI-J�k�zThKh�i��5צ�H%�$3H��_������׷�W�y~��i�.��3��O�m{���H������3��u]/S�|<\n���isʥ�}[��sĥ0��̈́�B�G�z�y�=�������5zij}C钪��%g}>~���Xه�L-#d��qc�zj��Z���-Ԗ��\�"�7�
�X�q� B@���2T�]g������n�u�b�:b���ǰm>�:r�J�Y�����Pj8��9��5���}�ө����.Er�'E9K+�f���鲾:MS|>��g�����d���{�ې�t�I��N�BY#��|1v�&~Nb��⻩6��:t����a�sVɋP����H�}A#�IY���X�*sW^��K���������:Yw�FGGk�I�`Ӻ�_�/��S������d�G��=KN��&h�f���2/Q�R$��i�7�3jqڱJmMe��j/mz�Kf�Pd��+E4��* ,��$��\�z��nu
1�V�R�,�$"�g礅*���DL�ԋ���]�ds�Z����%�Yg`jY��15+M�3aL<���u+�R��6�Ds6���5;Ӵ�X�Z)a �V�T�=�\�q��r����k$qp�{�'������ ��˕�
��9�ޕ��7��/� ^#pF����>�+��L��s�?��� ~P�D�����=~�o���N��L(�M1S������>��~���z�\F�7jq�#��� ����*�q�G۟����NS#L����N��9}>󭧔(�E8 �x�g��v��x�Ue�i/4I¬��(G�W�x?r	�m
N�il�f>��e<��������+�G�l�(Z2�k�6E�w+նS������|��kM��; �'x��w���}������ L���}����?oloJ/E���E�'DKQ�Zm�Z�:��<ȓ|\pK��?��>|JC/�o�{FI�\I�'ԣ��@�{���ץ<s��S��iqJ���{�<G!@�?��>�c�r]�����Y�C��}k7KӰt�������ꚽ��`�`�����ʐ�TkSfYɊ?mEcJ�0i� ��� �b��ª�{����֫j���_�̤�=�8a�O���\�>���v?P��{��>7�~��,�6���S�!�ޣ�?2:ow��;0�<��gR]Oֵ�5�t���L<L%��2�cj��ssG��k�g�h�^�UPUk�ΩfrI+Sȍ _�J��u���Z^J����O�����$�4�if�����t�:'�����|�3O���m�����?Pպ��:sB����]/C�|l�~��M����&�P�c�� ^�-A_K�$V�9����l��D2Gb�ܺ����p��xI���^J���������	2r�����Կ�n������n�j}7�k�=��WT˫Ꚇ���ƫ�OP��ejX�M����h&Xe>ʤ��w�f��=����L��?hR�!��<	�ߌʴ��#��^�_��<���?`G��z�k:���i0��N�N������q+T�ִ{Z)�fj�J�Qr@�qYԧO~i��jM_PVd��);[��a�B	�|�<J� ��=�q���r:�0�^@���$�0�;_���0�t����u\��gU{Ʀ��^�{��� Rx��ϯRv�5{i:?C��Ѹ�Z�D�ǩRVreS�ag��j��#��:��旦[�������h��B6�O�<��;ʍ\Ȍ)df�Q�鴨k_!.��,[,XHg�M����ꑡ�l�0�ȫ'l�H��GwRz��� ��{|�����^�t���7k{��������>��O�f��:7{���F��'@u��Ә��հ�e����L_�k\)z�/���v��� ��l%d��o]Z:l�MƊ�jM0�a�Ȗ��g嚽��<��ɻl��j}mӭk�u�;CYkF��i�g��i�±�Γ�-J�W�I-T�4�)vm�m�n��?�Y=������:��R�s�X+�>��5Һ���oI���gi8i�~���5
Q�N�����Jc�k��HPY6�Ut���:Y���� T_��M �}��_�	뮧�LƛlJ�Vմǎh&�rG#s�M��'�V�^�gwi�Z��Ԥ�j4+ ��&���{DK	c.�z9*O ��]�x�'�}����~�:���M�h�2s��O���>�cu.��Ұ��qt_izޭ���W+�K7/.�F�Uu���t� ���i��յ_x]ߴ�Tm�6hX���x���E��y~�3֊h{�%�ݏ��m�:�}gD��.w)�5
�+j<jU�/([V�#,_-4�N�d 
ٛ�������g�]՚O{�n��uw�M��^��tw�Orr�[�4�?� X����}���i}+�� N螝�����ãj���KUz�?@7n��*���-����;N�hb�`i�l8�݈ň�ޫtX�fnZ(�8�\ȺQ��:V�������=��ַf�K-A<�V>h��dt�F���\<����_l��G��g;��O������㽞��sO���S��k]5�<ikz�h�[T���ީl>�ԙ���k<���\�	1��xo]z��ꖝW��<:U�e�!�f%�"C�vxl��d��H�},���uw�#o��&mɲn���Zdv/T�Z噡�m>3<��~�J�"�����S�sS�?W�t�A����wm=�u?vt�c���jغ/'��U�����L�i�5'+�eAhE@A���?�!�g֢�V��]�[�!���i�� �!��� �95J��OZ�Ӄ@ַEN�ˡ0�x�)YR��s� z��B�nol�+��^�q� T�y��O}��tsz'���s8v�x�nV��ck]=�T��� �Wz�<1֍�ڵ�w���7j:J�_�������Xڧmsfi��<��Y8qa9�v��Zc�Tl�¯Dto�G�����G�5����f��V�ׯE4�O��Q���b�#�6�{@�}�{� ���W�:sٗL�J����s��>�t���vw���H��5<GAտF�к�]�Z�uHY3�m�X���]H�:Ɩ�u{��s�R��'MC��)!�FI�{�J��'��n�����Ӎ�B�X4���;�n�Eӭ�jhd�ØYO�	�HY��x�����W��u�GCJ엺L�kXX_�{i�^��|ƣ�A�6�3���]�m<.�p:~���[�6~�1SY���:s�܍B������D����� ���G�89�W��O])�i��ehG;QU�fV�(����yA>�`�,}/��I�w��a� �;ݯ�C]����ۯss�K]���a�w#Q�����~~OAW�NE��̴̔e��5�,v����oZg���}��Q�����m��-x)�I�	kUh��O�Y���MZ	bZ�Q�y��~�m�����=Y�5�ԍm5=�5�qMkPhg�/�H�j5Ů`�%�����G�<0�<)۟g=�o|]��=�{3�o��������gh�;Oc?��>����Q��Աӱ���OVVS9��ם�tG�}N��*��kf�[�o��nZ�Zg��r;<6���#2�����޳t���N��^Z�*j1�.�b:njB���|�e� .�d
B�y ��E���5��+�����=���9��*tEzé���j.Q"�֙ߝ���"����H��|�����G^7v��V�V�=C�z=�6�R֞"���e��~(u3�~�kF����	|�Ǎ���������ѫ׵�cD�g��e=��4�$�jpj��\�1Ú��{Zw�N��GD��������p��>�j�Ժ�zD�1�:c/�s�rf��ej�^6���j��qv���b���N�[E�+&��ƀ��l]����7�E��d��H�$������Ic�6u��b=��M����g��@�x)�d4�Ćg��K'�����z^��zN��gP��[�.����c��7��z��������������'I���f��ZcK*8�b/��I�6��Z[0Ʊ�!�NA����L�ye$��h�#�ݬ�1���.{���R�9�G��$��%I� �1Ǻ?n�:kF�{�ݎ�uWn�[�����/l�e��_��E�>YҺ_�{�����H6kb�n�eOWcXef�*z��Vhg_%��S�̪@���<{���$}�#/�d�I��v~�"�C� ���A�bw��s��j�/؎���}���˦v��?g���'3X��j�Z�Q���pmG4�vt� �88�PW-�-�4����8�~I���$�4��n <~��}�ӓ�7�����o�{Й���.����=t�m=?�._O�>�ԙ� k���,h:�T�������U+�|U/L�{��菩َ7�@�̤�	��
<�<� �>�����P����S�}���؏_���������^v#�uw���OQ�zN�l�ϧ4}�9����D~.#K剓qi��k0**%�uB��>u(U\��K�% �	BI�*��-B�5Y�,�O�R/�d_}�8?W! �ב���+ݾ��nOR������Og��� ��C���SX�5�;F讕�#x{�݋c�z�$�����چ��A������`���P�{x0�}Cq"�I���n2�>��ڋ�xf��qﻐ��(��j~�����T�-;s��uWi{g��Q��K������.6&6#w�tZ�Z&���l�hZ#GOJem�]JўH��5}BI��̒����h� �����I>��+��"Rj��>��X~��?ßӀH�}]�&+����W|�%	"��iG�q'�1bX���[�}~՚K|T��v�>�Ǯ_��ps��bi��y���l��2펔Ü�E�%ʙ(wm�?���/�|����������@�ǿ������)��=���� <�zv.��FF��U�B��!X�����y�q_����p6V���[�v��j��#���I?��}��Z�[
d��� +�~Ͽ��?8��4zb����\�5kŚV�P�۔�r���Wm�
����fy<�9 ����?���>��5#S-r�����{�_����Z����u\}<����R��eZ"������я�IQ�����	_r�� /���[[T����9o� rA���e�T��14�@���~��#�,x�gfU7I�!���YL��?�?$��jwgӦ��7Z�A�y�}�>�w?�ys�Vk$���H�����c�zȝ���R:�D���sRѴUԠq!���T�2�l|�tĤj�U%ei� ��\v9U���O�7��
��ū6�2B`�F�����(�ZN�ؿS�<~���ǭ;�RJ�WF�KrU�������~O�����:��>���+3��s�vG��!�ZoR�߫����]G�s��4�=�1:7�}�yx�[�]4u��=7S���eGC�9T6�m��̴�p����sH�y�'�LR���.��%w���Ի�]�Fǃn�ڮ�i/rjTd�H�F�O4#���U�� #u��f0����O���tF�y��H�����v�[�p�=����0;����v�2��k�=��y��߫��M}{W�4,]b2����t���de�f�����gh�cL�z��ٜ:�J�iڽkQO㥦�QBE����+-c��9KRGqG#�3nm�˯��w@�%�dm:du����H-]�&S�,XQZɒ?=H?,S+���/P{��E���{����������.�����kݸ��v;_��:�U{q�}�,���0�[6V�ĥ�gf�Uq�}5�衮��:�[��]n�V-�N��$��u��z�/,V��]�}8�>�l��oD�S_�P�F�a�8� {V�(�Zh߇�H�:7� �g�?[ջi�8�����WS{��׫��Ϡ}��Gr�w�^�v�ϔ4����ݡVѺw?Ol+��ظ�Q�0�H�0^/ԡ��Z�䆗M.��{jZ�WS�����������}H,��ޑ�ZCL�v�Q�</����ۻ{zi����(L�H���ص{��ĺܴ
�1ʝ��u������)��}����>��o�1�w�uXZfJ{;�U�.��~���k�v�9�Z�U��[˷�Y��A�0�\XG=+�;7bR�:<�֨�����$<ڡ�Lsj��u�~�Em(�^�`�Z�����7w�k�_Vb}�dZ���<ONH����a��I-����Zi"`a�c�L��3�$�~��&�����8��'�z�o]�}��{U\��E�E�};A�^�x�+���X�xDcb�o%	�y:�n5���,�.�"��XEsM���K O {��{�՛}
�����E��^(�;3N�>_�ߛ� <��#���� ��>d�������z��>�����7~����WG��T��	�5�s��b�j8О=(t׈|jQ새�[�w�������Ժ��4�3v��4���K�"�0��`<���UQ�%g����ޛ�u�},�:�����pS������<���H� ��HW���Wճ��_s}��� ��{���J�bv7����ޜ�����,J����Q�S��i�hƍ�C��azj'Ǝ��zŰ4����r��md���pV�7��m�����)4��z��o�d��	:������N���5�(�oz3Mm֬��̡bPd�)T�+FU�!;�햞����׮{��'އg��a���Y�t���&��ڧZ����Ұ:?���KFҧV��S�	��o�L\��I�e��n��t=GP����T�py[�DQ ��`�$�k����<�uC��t�zϤߡ�Z�!�[&*b�����g��:r�
	ٙ�V$� �~�=�{���w���+۟R��7���պ�Dj:�.��)�ڶEa���uf.>SK��<����6��͏�=����T7�/�t�:�W���rЙbP�*�I]}�;��2�� ��8q��x��x����=�-]���7f�4���ұV��xyVn�b�2FH���s}}���_��=��Ͻ���n~�:O�:� Ұ��N计��էK�4+�E������uf8�:<NJ	1��� �OL��K����H�]{k�Ɩ�D�q�)w#�ia��gAد�%IG"���������e��L�7T��-@�Z�$ԥ�g�<�p�\�Bd(9���1���oZC�_���3���cz��x���ڎ��mo�;�Q���O�:�mMrm�;bgd4�N@���\P�i򿥟� ^�_�:&�%r��)�k���fk�A^����g�FU=�\�OMz����{d�]gJ�V�
9�Bikv�'5��5���ݢ,1��:�+�����'�n����?����;o�n��ַ�����}3�X����g��V�FFnV�dd�Ac�7dui�U�>�oOv�J��e�V��|U泤��O'���E��G{2:�h��׸g1���������N�*�����b���ijJ�!k�"N��,���evH��k1���k:���Ɵ�}��A��PdNN����O�^o�y�uX��Ff����IYn�y����F�]E�`k�7>�/s*ئ�����he�' �3֔���(�v���z��m5�:mT��/R��Ѵ~�J�D��#��؋�g��J9#���=�KG����� O�뤙f�?Nt(ԏqr�,FNV��,����ZRg��m��"���l�-�6��mQ|Q�<H�x� O��<G���������X�RD�K���Tr�� ���܏�� ��>�����N�v�ۿn��E�_At�������C�OT�ueGL�o����i�#����7Jx�q\�ޥ�'6�XC'`+8�¢�*�F�~�*����f=z/�ú�G%���~x �E�h��~ٹ���S�{J���{d���.���[��Нk�]��NCt �>���,��Q�ؕ��n��9^\�'D��Lɸ�έ���5z�<��h�b�����-����=+s s�9sȑ~�%��7�����xPO��щiY�����,,z��Ȧ=�-� W˱X��O
�E�X0�enET5�KR>Ge����������@��OJ#��g��%�>Gv���
�#`�ı��G�� Yw� �b2�xyvfT����C%�\����&y���d��f� x^�{�?j߈�
�cF��;(��1����*"�"B�t#'$�D����-�����r����:�	c���R���SB�OiS�]Դ/BӚ�FHK1�/(l�M1_�)�Y�?"������Q@�5?�T�* Ɣ�Y��
,���2�L��+�j�&
��gc�0��Tc��F�u�Ε_�|�<@*��1S������;c(^s���*�o�Ԛ3m�l���y�� &H�kR�Q;�l�m��r��쿓P�X�%"Y���c:�f�k�)�7�,��ʭ�[wۓ�� �@ 1����Vɒ���Lhe�I�/�Ȅ-A�qݚ_$LlKzcPU�ŉjH3�։�YBDR�dnPq�����b�B?��c6��3)J/�#��2P�Iq��V ����X�hUk������I�w7�W���� oLd�JR��,�����.t�#�^*AEUB�r�v1��/���ҝ/
xRiO��hː8�ј��� ���F�a<k>�CF�fY�Q��6(���-�˷ߚ�crY�9cP���-�iT�ʭ�EU����U�c���Q��2�����vW��;2Abľ�0������-7b2y����"�c+ϑ���з���(][���:~E�;�r唆��ߊ��Lel�;*���R<�%��� !���c��`���<�5�?�Ɋ&ƕx
Xm㌜��ll{�G��nŜ_9�x~��[&�z3y��[���Y�o��=�m�F1�H	���G٭J�,|��~Cr�B�6�G�UcU��I�Hbc�g}Ӑ�+�dO�b�	�RY�O�\^"m� |sVx8�5�A�+.,�e�c쌪�D5	eIz��ג�%��2����X�,b8I���I�84��2�y���rŘBV�d-����X���yG�8�tTt�T"-Wu�-[c`�#�J��Q��NS�2���U�U���DD+L�4W����!�#e9bDqv$���"�� �ձ� � �  ��1�����]��T.��CL��d��v�Y�U%�� ��c**�FP>vM��&�F\�|�f!Q@.8��>��h�9ɮ<��%�h�XAV��$ޮ ��� @�Sb���D�y]��q_�(̂�(�FR7o���=�:)�sFzQR��QR��n�S?��#�PO?V27:~s�6�F���W+��t���ۈ�!��I�錹s(!T�Ntl5{�+ʸ֭��3B6�By}Y�1�R�5���<�SFp�~;�F��UK7Ϧ1%�WZ-� &�f|�?��&����r���J|���12ɚ*��VƱ��f>9Bj�|���8�[}���p��kfR�z$J��_�d8�8N�K
�bX�(�V1x��,))MN=�d�poM����Z��ڰ�y#�6SPӗ'Yd�*Rm^l��`�fU<e�cR���Sa���|ʥ����
�E���h�q�I���S��<`�h�oƴ򞮩�6���/-� �͵6%�c+.N��Le�����Dц&B��UN�Vc�����).��f�^(��q���/}�nID����v%ޛ�������o-��Ƨ�R��L����<0�	d�.�i������/c��oLf��[�_At�:cj��8d.1�d>C4��M2��+�?�E���D��qt���_oޏR�5)����Đ�R@ ����/ }+/��.��4-զM�n=&kK���lFA �rO��2H9��;!��3�:5'����p��"	����d|�fS�i�eQ������,jUX�7�z�n�d� ��b-'s!Q̎!�u���Ge;G9
�vo�X�ё��ڟ�N,�ƭ>���,�ƆƥAKp÷��B�hI�^�Ѣ���o~d��v�{ï���چ��3_�/�L�����e�U��`�Ӆ�ԉ���vǤ�c�=8їJ�5g�4�8�a��<I誣�� �C�#�joZ:=�����]�w�iڦ������<�pU�DN8�9焔�Aݝ�ޟ�_u}��{��ο�/���vcK�:S�4���ZGQ���C�:_'#�5JW�6�|opkl�)%�s׬�	��W���C��滸4飵4���%(�b̵��f����D��k�����IP�>�|J/@�sWf��CӴ*��X��+-MO媥x�ұ.R#BK.��`9�G����'g��7�O�R{9�?q#��Z��� u{�ޣ��tOMSH����Դ�����l�[L��i�FvO'*��]��d�����Ӻ��7�7�͝5��t��f�Ƨu&��i?%����Dh��,ʨ{�?�^�o��k�:U���Ϩ�zU��]�R=h�e�o=K���y�A^9gQ�;�Q�#�����?C�F���>����Ϩ;�0����a��:�xW���ӵy����4��Ȣ�pmA9�N8A�o�� �/e����v���ý`ժKx ˊ�1�B�l���#G�����z����U��,�<�x=�I7�y�?'��0+���Ӟ����;�����@�wxp{��BK�=��k�#�X��i8x?�t�[QǎV���iZ�YP�\Id����F�'������(u����Я���D��`�v�#W��[G*!�ZN��ic���{��f���un�Ž�:�5E�x-ӭ� N��IjJ��*	"��ч��A�u�Μ��Қ����h�SP�m��a�=��x���A���KGBү�꘺�.������A1ĝ22c������_�}A�Ƶ6�e塧�f"}R�R4�l,*q��p�G!<�deU4���7q|S��q����Y��޽uR?��Rey��8|�y��#��8��Ch?����q��-�#ׯ�|/����w�a��P�:��O]/I�s1����t��-e� ������J��X5�TA��Z%�RH8Z��nX H.2�&�� ��{�A_y�Z��Ht�ګ�qLP�ҡ�|`/&Y(i�E�G�2��ל��o�ݽ�`�~�� �O�.��Oҽ��\��w�z�X��[�������V���Yb-�1H�Bќ%�1c��||(���B���卧�رam�*��/w�Yk�v�1�$��j���>�����g�έ7M,I��c����Z�&�,�IV9��+0�A/�8і9�x�y��lg����{��Oӫ�a���� q�ֽ��9�Z�^���KB]>z�N��Z���|�r��HV�k��-����W��_]9�F����[�wj�э:�_��5��)�Yf�C
����G!h�g���[��p�Oh��55�&MF㸳e4��6`�pׂ�:�ʈ�'���ci9�=���ҿڷ{tN��'w}�a�[�\��W��&&Omz��t�bn����t�K�:F�������$!�=j&���� lV� �ڍ}3P��24ˤ��Ǚ�"xn�~v�v�vQ�?jr3n����~�U�q�)f��N%i_�̑�*"��*Pn�>��$��x��2�������r}��^��=c��?h������~�����^�͆������-N��4mM_+T��4L�W}5�l琾n�{{퍿Ց;[��j��{2��Tfjo"�`�Nhf���jG0e�7���tͧ�����EkۏE���h U�eג�Y�
��Z���~^�sJDS9�>8���Khzl5N�����u^���Ph���+Eִ-jqJ�U�
�i�zU��L|��:UC^�Ș�?�G�Am��\B�3v�wI#?�fF �)�(�>NO�>�f�O^�RF���r����#��{���3e��.��6���녔2r����H�>���r��_%���d*G)qݗ�RS�����e��+�_$�䏫��9Q�?�O�>liv�x�Crx�<���rG�g=�6�����Y�ee"��a��d���1��Ic��w�jRjZ�y�9�6 �{@S�������V�'���O<�G������ۼ�.����v��)a����4(C�E��՝��4�(1r�V;bSպ�i%�#�9ջ��� 8!��r��G���i5��>�w�y�9�u�O�'���}��' �] W]�o�҆�حI.C�m?� ���'GRY�%Q�>�jZ|���g=����� ����e����;���c������y�=��a��������:O�z�Xa����S���<��t� z�����]O��h=/�xZB�١�e���)H�[���]�o�MJ�ˠR�
�LL� 4� ��Ռ�ۑ�v� ���x<b/�JS����c��Kګ�'���t�<������ݛ�ޣ�\�ܯ��� S��h}S�h=��~��[X��t����:�{�9Yz�lz�P�\����M�c��Pl�e�[6P�v����Cgu>��<�T��C�#G�)ORêL��:3����L�B���oU�M�SbjP���Y�U���7o�b�|R����߯�H�
Ȭ��/�_�߹��v㼞�����h��ugK�aӝ��h�!�'/K|�����S�֪۠uFļp���9�����3$f��6�H���4��Yv�b:��q�ivg�E��M�Pp~�,݅����3�+Y����[{Rگ�p֒W��	Q��!��X�m<)�&�G�ȏ�v@�?]��;�jtN�vW�gP{V���t>�{D��f��=���i����WOw+��66��K���5�W''*�5��r�gm>6z�НB������_[���nN�/�_�j�fHm�{��f$ET=�ys8^�u���o]҅x��6F�i��JZ3TD�ğĖ������s������u��k�s�{B꼎�K�����,m�������zG�)x�q���e������"��H���Y8���������X���-ú5�:v�Ӎ�'�iۚ���~iF�j��.�������7���V	���Ga�n*76�PtU����F�$Տ�h�ے�y�x�(��9��:���;t� ۏ�sڮ��oc5n�f�����k�v�L�-kO����i���+��c'�u�#U��� C�Lq0��R�t]3�3:�Xx0��<{�cd�[M�6����p[�A��W�z�#X��=��S�W�-�����>vRk|�6;g\��u�khpA%�Ni~f�4�+Z����R���#z�W�f@�&�1�ߟ��n_�.��t�Is2���ڶ��]Uٛ�g����˹:�Q�v&�ݮ^�J]��(eKM�P�Z�k���1_.���=�h�э"�Y��)�[�j�Q?�Ε41�?N��k2���i�S�!��K~7TN�����i:�pHGmzsVH�i�궤���]����I	B�>zަ��`z�_�}�ϲ���z+&y�l}{���ޅꃙ=O\N���޳���������'�-���J׭��)�n���.��� � �z̛[\澧�U�VM_O��'�pifH`�;TE��)�ڍb��f��v�:���A���/�>�䋙��ᬍS��k�3��Ɠ$�iZ�Z���Z� �	�{�]����Ӟ�u��v����l�K���٧i��V�.��5.���ߜ���^6�M���9:��b�j:�t�TJ�t{m�ooj�`ڗ5�gI�j���z�R�[��"�n�ܰ���#��m��R�E̊�V궻�}f�������i$�M"��i#���� �m�^�X�o��)�B���#��=�~�����gj}�u����=��s�;���nߤ�'�}�:6\:oS�n��WWŎHi��剓�=3+�����3��s�lo�۵��_e�Ҵ����IM*ƣ%�iwU{KnS+)+GD�4Q"�̡����ݦT���{SE
5zm�-D$��֊�U��.�(��(+�+0�x�q[�?�k���#�W��wtzsK�� n;a�S�!�:.>����0�����Σ���gs���r�)1������h}4�� �n�]���&��z���mi���C�^TiQ$f	@��!�34]�tKpo�|݇�eն�������U&W��m�x߽��єI�5w���;�����׺]��;�o@엲/o]��:dw�=���N�^��t�+�5
�Y�ɶORdfi�@�:5�.U<G#�#5������|-��{��c@�u�=���j3�V+2�h�"4U'�3M'�X�7��c�1�����6��6^��c�4��?�Z��0y!X��x;��GB�'�<j��fGR�s�q���E�G���%���y�۞�j���:��{������:�A���n��.�}Nw���3����3ed��a\ֹ���={qXQ��*uibaV*u�������G���̏�v&k(�ZD��7��O���H�,�ҫ�K1�qd�h���l� p��1��Lٯx}K��c�WGн��Q�;н���_s�N��-C����c�N��.�v\����K�?�U�e���ӳ��j�L��ޗP��%���T6�;��ֵ����X,�%��;k�h"񷒭����H�)j��sC:���~��U��r�z[�;2MQdI���#*W�;3J�*�-f��XdB,�
�9�{����K�݋���3��B{l�7\�&SvOD�N��o\�jg<:g�z[K]��Ȍ1�^@�6Vt�Pӥu���!�?H�/��V����3n��J{W���)�m�+�)���9�b��"����N��M�����0mm�v����;14�4� ����<rH�4a�\�� t=� �O�^�j~��Q�P�� ����:O�4}�{O���V��;Z�qu�t~�9����&x��5���(2���)Ǐ����Pu�;S�o��2Ĩ!mN�S�l�R�_�Z:�+��7I�eN��z��� �.�Pt�Ԣ�Z�1��R����<W^�{3ʥ9��KP��z�O��C�ӧ��u����o'�>�:��'n��N��-c��	\-?E�ÏYtκ��{���fjy�}t�n)�,��K���#���u�nnMxЋti�m��O��,��m$2�E�f��TWi�?��Ś��<���OG��ֶU�е}m�ײ�L�,AQ�X�x5kp���d��f���9��~����N�:����W�}�h�K�<��o#�Gpq23i�#^�h�D5M7��N-�g|���ez�7~���D"��ؕ�ꪇ�~�.�3'���$�FQ}:�G<��H>����ٽi�ZVm�n���Vg��ӛP�_��)İ���L����HZ�}��U������O���^�vc������ ��M�R�uҚ�MS�y�]W�rpr�λ��Im�j�ǖ��V���-�{v�s�-N�����d�e/��{"�  �A�܂0x9�zm]nT�������aGEZ%Dg�;�N{{��@��?��ʰ9������v�GFl���WHv����޸L8��V�5Θ�Ŷ����m��Yr�nV��y�c�*M
ڂU�j�P#��X�a`x�&`	#Ȝ��t����fPW�2{X#����xI8�G�x$s���ۯ�k���}C����CZώVdt������&�tn�a�ޮ���T6E�>�o!�o�V���׃��&X��=�R����g�kd��1x��#�'��>��=q�z���a�}�쇹��?�=Q�~��:�N�UL�����ƩL>��Vプ�^�������i�;�Mä#,h����IbD�$=�� {'�}�������Rˑ§��~>� �׳�w��WH�>��۝oU�u��?����=��6��u�PWX�|�|>�Z&_Gtmt�Q!��hd��j˵���ݝ!�dL�-�"����E�Ȟ�N�	R��	�X��bkVj�H�ǆ
�I��o��z���0����?s�����������3��y���-Uղ��_7,��v4���gP�1�]RVt�e��c6J��.�?̤F+���(xL��G�n�r�U4mA��ʕ c<� fU�?D�W�׎3Z'�9���~���x�]����U�r��v���|��׵ uhg{��ލ�O�����5����k�Ϗ�jXjO*�ܚ���m]!-���RC�#a���!y��zET�%gG<�������%A�A�9��~����S���Q[_�R�����:7Lt~��y��Ct���:vd \lY�Ч�*�K66�'y���}�}����~�O���#헷�����������}���nڌtȬ��/5�g`�T��a�������W.����|���x� _��sq��;;���q������m��b� 0�>�s�*C��@���c�����?g�Ӥ�W�r��� �KF�Te�W#�������}0<o
dHW�_�eM�5���-���$�N��׵">�F��~�=3����?�{�2����o����C���� �_t-/X����~&6N5c���D�v��eR�n~7;�@�r��-V�Uh�DÒ�@=���������i��UW)��$q��!�� �e-A� N,���6yt���|h��+�[��I�V��Pl�G�l6��tڕb��j^HG �$r�z�߯�q���%X;©>���@�O#�:N�L:h�ޫ�Fyt���K%��i����$\)p;���T׵eI&[�V���,`����O�O����i�hh�j�<�w]�>�� w��wC/��} 4@˿����:�@�:�!���Uצ5'�wL�}C�M)2�ώ=�1r��L?,'|U52_K6��Kr��p�j���,r9<��;��B}D�"�r��X���B(,Q���e�2�~�?x��n�X�J��/c;�l>��s���n��/G�ët>�u�b�i�^�{��F:~�՝K��'3D��i:%�":��#�FE[&�^���6�n�-��X,��fT�_P�x+��iz�ʬc�v�֓=��[�'?��@ �Z��Է��v�b��k��򰰾�g�
�������_�`{-W�3�����߯o�����g�� B��F�^��wc�}��}�� ��W�z� Qj��T���;P�Vn��hS5�E�x�o5�.��M�{Z��o��ojl�:zݿ�ԡ���Q�]������)�� 3�T��m}���ޫ�hE�{�R��'���Ջ
�M<��ġQ=�D1����~�{��5����:��힥�~�kV���m�oJbi�9z�~:�
������S��zv��W+>�I]V����G�V��{���V5�����덽��M�v-A�	�"�����+�ig�K�X��b�PF���o���h�zp��n�F��ӯ$:m�=#.��H$1�$����R�9�>���k�OR�N�>�.��Ϲz�v���w�����v����9�n��{��1:�S��\���S'2h��F�M�{��n�j[ΥK[Ҟ���z��='O�(i:�������xV�2�3Ү��Y">�X��U��I.��[ڵ���l۷wK�/�h4�q�)�X�ʎB�:q�J=�����'BvS��I]'I�O�^��=?����:�t�w�{���2��s����3p�0�?'*''�:y��x��%��s�{W~����յZ�R�3|�������
!B|�W� �2��s��Hz(z1��z��u��<�TI5� S�>�2�AkfN��'4n1�K-����U��&�������� �˪�5Mw�})�iv�=[��#M��#�5L�=JGGY�i�s��q�2&��7��g��kU�c\����?κ���;�T0��$6;͚���:��pA��D���B��S��rU�:DIޢ�<R��%��H9<��}����Nbu3v� �V�$Y�]���'q��̓����w��1 �+��5���?"�:�}���K�/M�]A�G�hW$b���碖T���UH>���R��!���%�����gսwO����Vh��K�]��Y~�ǵ")�n�%����]c�Wz;�}���B�6��ݺ��+��&�Mӝ��n��y:M2�.�Ыm&�����.8tȶE5�:7����z� �o���'����<�jd��rCe���V�0I���#ZӉ+����@�v��{�/Rٵ��t⭫�Q�E�b)��*V�b+,����-y"��^)!ή��}O����헷�t=Y�=����u�nrt���.����r(q�Λ���S���Y�#Qɲ	&B��zۯ�=��M'pC���6��t�WF�vn�Ԧ���8�O�֖�O�3�)
+��׭[��:֏kil��?�jv�#O�y��f7_�����y����4�"������o������m=�wVZ4�pL��Ja�NCUmFG�Ϗ�|m�)���/~�=F��,���rI�h�+���� ͚� �e�ؓ�H	1	j���u|�~���"�� g�޼Ox��5�m��{;퓬{e�,��wg�g{��S��vT�iz���z���_N���:b�&��Rߏ���8��m���>���m�,�]��ڞ�ޡ$��qڲl�c�k$�J�0��NcE�]�YH����WC���GI�P��7>�J�Rث����Ek� ����(��V#WVU�����t��� ��k�;�����������S��e�9}�� D�&��RI���$��3F4�Y�Һţ:t��p�7�'V�^��u����i�jmB����g��Z~I��%�˴r�#�R>��I��[�����Z�=8�__׷�ԥGMH�8������g�
��4h���P���9�_�����|���{[��;���9��n��.��z�M\=��\>���&8ea\�����O��K�wЈ��w��X!�4�W��Ƭb����x�����g��\�C��U�U�T���B$��_���=�p}�w�����>���������o�����ʖ��I�g�����L}' �m��l�.R��V��hN�T�&:���՝st�Z��ô�P�r�I�WZ��I ��ε[�f���g�ĮB�Tz+r�ޙh�g[�SG�qУN�A�;WJ �s'��¬Oeb�H
�ȣ��#׽�u�n���S���ް�:�O�.��^�������Y���z~?O�gTi��1�t0�<��o���S�m��z�)�,1*"F����i��<2���-���>��u�eWD�rŞiQ�>ï=�ܓ����~73�Ϻ�鮃��:�Lѽ�iZ�`u�����ah����A�>�ƅ�=_���70�y�jM�ƭ	aL>B~���X�����q�"����(Ѓ��V@O
���M>K�Eb�����	Y>���2?��x��9E��8���s:K��A�{m��u��w_��CJ����_zt� ������st,�o�]B�lt��YQ�hڥ��\�x�z���BU��odr�>�����s��;e�Y'���\�/I��������?��ݽg��>}�����~�=��]��o��@���i��k�w��4����h��9j�F�+d��mkQ�Fћ���������@���fx ���˞���9�a����L���A,��x�~}׹]#�[[�'r5\�^����tGN�a���K�gi�X�Z���Q���=z�K5��8�\�LF��Y���J�<QW�ـ����pH ����'�b�����x����)?O�=�x��|�� �n;s��w�ڎ�]���x����c��z� Mi�-�l=^^A�cO��kc�X���9�u��cJ�'��F�H���G�S�<�����	�/�uz��x���	���p������c������#��#��>��J��~�����ږ��.����O�jk2ui�89P5
��x�C�͂H�&�{[�x�D=�G؏ϯ���U`Ðyo��Dk9r����+c1[����R��s!T����3��2����R�qF���a��pF׏�#���q*��`���R��T� ��gL����㏔)�i;�λ�Q&T��1OA�c[��� ��W��D���Ĭ�YA}�� c�'[**�:J��[���(��6�ǀ.��Y�~;1�+M�,�WȲq�	�~)ϛL��!G��o"�g�n�x�$�L�қ:�GLY�����i�K|�B���ı�琲[�I�ӕ�`^��vw�<~
���vc7/��u�[%Vĺ4x�9*��uBH#�RX�DI��{�J���5�j���ZO!p��\��¥f&6@�L�3_-@�V�j�#0�d��⪭��+ � }����f�0��ϑ�bNu`���5`*6*?y�W��cڇ����9�U&E9�鎎|���6�l
rA������x����X�0�����|R|�.*�Fc*X舨*�4����g��˚H�h\��M[�/�1j����rl��:�oܝy�i0��
�'�C�� :�EY1���ќ���&3�B�3����>E�|��c�Ru�{Z�_I��yO*2��`x��R��.�Y5("��Ł�?�[3�j�
~`f���F�S�v1��U���:W6f�*@$~��P£��K���7�H�~U� j�\t�c�`�y��0U91�"���E�(ҕ*�i���*����+q�
E�����s���&�~Y�ʕ�Ì�IY+Tx�Hf��� B����8|b2����L�V�BP$�X9,�?�� J�6�cp�])98J�%�=2
�6C�gU+5<����c�h�:��
��[Y�t�Fʰ����+G�Vb	��a�=\m�\.��/^�ܼ� �4��ˋ�O�1��K�����n �Fftc·f�6,� .⧊�;+N�]�~�Ce|c$/AC4-5f,�0�j��.Wf$1�����r�S�3��$�l�q��� �Fw~L�*��XŔ��_ vF�ŉ�@��#��IR`=M$x� l�cJ�5���Q��$a%,J��������f�_�]�m��b�R;�� /��H�.��1�d���S
{ҫ��˳�Y�Q�n,���6--C��Nn|���t%RLmV`c�m����MǦ23����:��)��)���M�(?�N��]��7 E�NN���Q� Q���� �]���͙8�%���c%9�D��d��-[~<k&�-Ul~�/��H� �7�[����Lx�8�� ���<-B���(y�r6hdd� ��e�Q�x��i+*�#��w�{���c3���˻��~�Nw���\��dZ!qQ&٦�@��e���;	cU�(�᷉h?t5P���Q�
�pYW�
�Ld���	�R�Ǝ�9	"9����%Ô�P����JMj��N\<X�ӥ�kZb.-P�8��z�e@���2@�5g��ˏ�r dx�P���.<�e��9ԖJ7��D�P�"1g�6&;�E��\�L����>uf}��;��6c�FG�>)R��<ъ��������Uٸ*NE��p��E��	�1/�8����;�ѳa�r��Q�l]�R��c<7S�ĵ�qH��N��I�1��V��Mi>/*.��BʜvQ���vNڼ3���=����'�ixo��{�~6>E&+��QTJ��qʪN��c9�֝��zv���l�WzbW"T�EFpȼ����M�X�8d�چ�1���:�f��%�! 4E�t
�䖗�q�� �K� }��}���������W�u5����\��z�nQƄ���^�����TY��/8�A�gv+#�n��Z-e�u��;i�_���g�㺕���'�W�d��=Ą���wt�J�_ph�N������4VJ�Bj59X��Φ+����q��^�~�^����B�zTS@�,�:��=X0� ����cJO����B�eɀ��yƟ���Wըk�vlmLZ��3�DLW*�G�r�%�{ �����%��\k�:Əj���N��_Rd��ͧ]�ҸT$r�,<b��8���{G���{y��12�z�����C�:X�-��/�3�k�c'7T�v���t�}�r��{�b�#��|/)q�:�g��q�w�V�hv>���(��xko�VZrW�䮆�q�ᶋ,����ou0�Gv�R�;�c��=�>��:Q�� �Oo�HTن���V�|�YI FxdXR�4��(���������gNuGX{���M{��� v��h�_�{z����Mft��I�\-#'R�~��֒�����d»(�i�����M����Ӿk�R��O�_�t���*�mP��O$lZ%�)� +�Ѣ𻣨|xU���>��s���z�%�`Zzݸ���*Իe�)���,�!'�6i#�{��'�>�����@��t���9:~�ѽ4�u7U�t���X=+�>&NN9�ƞ�YG3+�H�Ra�:�V��e�υ�J�N�X�	ۭ4j튱\�ey.�^Ri�(��3��W�G���m|.u/�q\��m���5ަ�N���:B�RK�,=xk����Ei$gvx�baH��㫿K���i���� ��o7�� Ӯ�h����:��_]�Ӄ���9���Ȇ�4��L�;dL��W��_Z:w�'J7V����e�J�J�j��^�j�b`�]�G-i~�b�Q,r���]ߟ	ڌ�M����;n0����Wj�N�jh���X��$H�-gI�$� I���I������ Z�w����z�7�y�7M��p��v����N�%Ԙ��r:�cY���$1H�Vb�?�IOkj�4;�)tj6c�Z9>fɫ�c��cp#RDIf�S��_�D��I��â5[;n�Ԟ"��S��y��k)�YX�X����ؓ�����l;����������o���\MG�}��MSU����Ӵ䶉���]/R�t�i:s��9!�X~FU2�)����d|)��/����E�؞��%�5�Ѱ���c�	ȃ�+�m(X!��;�˦�{��ڦ�y%�T�U���|�ԫONp�-f��$�M{��@�I',Q+�}����ݲ������ Zk�����^�v�=:!����v���s�%���Ю���\�Βș/��<�u�|�����Ӿ�i4����gZu�ik=I��J{���;�ct��Y𥗾9`v&��� 6:�7���.h�dU�Q�K�Cv��	��$�(���d%%,$�*�f�k=���t=k�~�t?`^�;;�vo�ս��[�Zާ�t_l5\�juN��t�$������ҫ����ϕ]����3�wFu�6֛�]����X�ze*�;S����%��U<���Z�q��t���}[�u-JqT��t���$�^"ݦ%��&(���
�Y@\����{�� L>���?Z�5���y���-н�պW���~N����S��nL����wk�Jj�x�>�1�
�ddjy�C]a���Դ>���oI��ҒI$��k���ey��\���k�/l �/I4�G{~��J��&q6�cX�4���Y"G��{���I��|��>%��&�9���PuK�*fY�Ͷ��G��іJ��������Q<�z��\�Xѿxܶ�
1E�JZ��nCY�\������k
��٧ȥI�]P~��S��W�y��WZ����Z�Y`�bGR��Z�v���.�:n'<��TţI�&�ɥ��v9y�S�in� �/${b�Y��;�qϥoA@񘜺�i1��iO�x�� ?�r���؜�N��tΜ�oK�^��mT�f��u+�ckL�Y?�L	Ә�όn��ŕ���N��If�kr�h��G����rG*����e�P�p��6<�T<�{�W�z�	�� \}���ѝ���=;n���櫚U�����s�/~��iS��e�یr��W�x�Jq �ܗkhv��$��i�� dr{y��}/ܟ]�,�ތ���)�5��yP�C� �,g��}\�?<�/���O�����>��7wz��N���Z�����4��=�{��BMF�����~�Ğ��j����x�Pix��N���Һ�C�i�o�uQ�ݧi�	-���G��H����Z	�$d�,t��y�P:����K�kV�o[�$qV�W�#��$�J�WD�)dX�Ê�,��<��D���G�G�ޤ�O��ڷ��{����e�S�wcm}[�1�1���g�w�|z�+�u��\���s�Ip����;Sf��>�l�N��ݕ���x�Z��7s����i��x[��D1��rG���V�.m/C�C�`x[�D9� k�jB�b���d�T/ˢ��i���'N~����;��C����}�uN� E�Oz]�l������&N����;K�kZ~'\�Jt�Q�ErcO���<*�5ӫ�;�v��T��]��ُɶ��_�ʕ1.���41U�9��Pv�&>;2$���>���n�{a�_T�nC1��Xy|b9G+h���b{P��?n(���.����j��~�����޽�l��֯���������l=��5�.��j]�ӆ���az�#Ϗ<~���MS�������i����~':��zΤ�t�S�ڤu� ni�]%�It[	"V����Vm:y������*{�f��Z/Pz���q,Ri��I�Rx�
Vר��5X^-Z�_td�QP���q���l�����{����������.��u.��W�=M�5�[O�z��n�֡���i��>�L�[2l"��'�.�.��gU�̕*+%�"�Q�\�,JʱM�ۭ�bF_�vx?���=�[��WE�(��?�y�j֒�e���g�v��%�*D�l�G�bc�ts�^�}��y���b}�u_�.���{����CD��i'X���oC�o���:������#�qo{�]&M���>�{���۫��i���6,U�*n�嶗5�����d�R
�G�*�������C�n�R��v)i��am�-k�я��u�#V4#���U�<�#x��'f]�����4�/w]I�^���v������v��pzK�f�Қ�;i~�;O������|l�d���i]S�N���P��=c�?Pvo�uMG���������m�~��Wu*���k�Z�ڟR�K]��%�Js����E�[�pZ�{PڬY�=��:~�:�o�g�-=Ǧ*�+��#�
,6]�Ť{[�ً���E��}��j�̌��{����i�#�a�c����:J�����μ��N���u
q��,ō�߄��n�U�&৸c�:�m6�Kjҗ,#��׷%�0S�m��C��Ǚ͏���4�kF�4m_n4l�5� ڦ:����3J=B��є=i�����s�r{���{5����N�u�ip;��鞏��;m��{��GN���ҴΉ���Y�ˇ��҉i��0�&��F,�P��\\�Ɩ���Q��Ε�[z[�mf:5��K�ze[S˨-S�z�F�5��X4���^�����ڗ]���/Z����j�"�rJU�5TR6D�I�-��H�b���֞Yc~s���=��'Mu������ zs;��C#��uн���(uޟ�ѵ��c#[m>0������}-��M[RD�6C��w����5^��gh�z����[J3i�[�j�`���3��	|f�H���6��\������;�bk�������1ٱ^�k�Q� d�6�V��ȍ�b�$,0�U���=U�k�����%#�ۻ��Ku>���;x��P�,�@�`k�0����Z�Ueʫ*� ���ދi�ݍF���W�l�Қa���-��=�2y�j�M��,I1=���=m�w��^(����~��˺��,v�~�h;F������s=�b�����Tw������7���?k�t���`�[��'.�vV8Ѵ��K�k,_�Č��L��͖=������cO��J��۵ e2Z1���nMP]�N�#�<UUI�^I;D5�D�(t+���)$��w����a �e5�էFɭ�en%,��ƅB�3Ywy����������Bwǩ}�v߹]��W��a�+���u|���մ��2�=_���\܌ތ�
� �)J����:�iZ�)c�0��.��W��.����S�*]�U���?��H#�+����SD��;cx��7��eVKzM
��r7�Rޟn�s�n�,���I�h�	�<N�q�D�|gU5Oի�7Qh����^�헽=e�Zd�Q�ޱ�F��q�f�����:~���S����M�p�ϝ��*�Cp��0�_���=ô�����uj��KJ�;Q/OU�U��T����+٘�sPi|U�v��N���ժ��"��X�Os�U�CF���i!�O�<������h�n���>��W����Flݿ��W2���z~���.�^�Һs��td�-��_#N��Qp�/��W��[��+գ�Θi��v�%Id����ݵ�	ϖ}F�v�Z�&�7�[+��'/���U���nn������ߚ�H���եZ�1Nb�B�9f��^88�1������~�ܟi�O���ĺw�wn:N�]�u�CC#� J�Vӳty�����6���7$	�&���{����ϊΡnN-E�����-c��%��<9G�+��H� ��=�JǖI��sf�����M|�^�*kLk��t'��;�Ɋ2�H���)�t�(dbi�H��~�5ޛ�E�'�����#�b`�㺚7F�_Sdi:_�u��|��S��x�T��&��S5aב���Ю���Ӿ�=j�b��.�Ri�E]�
H��E(Zܱ�i4��3��� �,t^��r̲mM��l��Y �B�U��}����4�0E*_`ʞ����5���t�l�GUu_04�s��:�5�� ���7]꽦�A��I�����?lr,jn�i���x��&�?&����.�׼��_F$�e��Id�z��b{�Ee�` A+��Ay��m7K:En��z��E�:��2x��[�镕Gd1� 5|�坌Hb�>�ݵC����]��Oa����N��}����_A��΅�����h=f0�M'P|�S�L���㾣�5��r�ƋѬu�ޒ�]�+�>���Wbd�'�Rr�|��p��S =�z����ZĮ$�f�)��=�6����ó�!�v? ����-��ϗv��ߢt_��^�'�/�z�24�:���%������ca�_�J�rsc���jc�&����*Fݿ��ݫF Is�<@���y�T�j�4d�K)x'�{�t � q��[��}}�GZв��s�������l�n��\�G{5I�bj=��lu�r�9Tt΂�Ӽ�+S�NsX����^J��+ϿC�>���=s�������>���x�Nd>�~�zN�]	��:�S��n���N�{�f�n��zN���]g��Yvã��¥�\�_1��e��t�Z�����V�w���������?<~	�r�t��+�'���?c������_Q��Zt�;#�kM���E�WOv���gL�mS��=/����qzs/YeW��1��y��8�DM�$h�1H�*L��q��"�  }��C�S�<S� w����z`P����;����i��}���UuMc�=���i�:Oqz�=[���ٞ�Ѵ�aiڿ[�Xױ��c��KN��q���Z�t�|ɧ�_TwV�5	�H�p�������U^�`
�;�g�m�ݗ`���{<�zn��!'�LIW����3�w'���~���o�9�vE�24��5Ԛzi=��],��^�ھ�Gx���h��K%�����N���-Qj���E�M�� �"�$� ��<39���2���^�q�}~�c�M� ���B�@�~��O���R�ȥ��vɵ2/ZѼ��ɽ�E����h��KϪef�;9�{?�?�ʣ�1?n?��,����Z��1jx�q 0Ur
�-��v!�� �Uq�-�7 � /���� �g�[�߿�� �z9i�6w�?*ت�3ƊҔ�Ģ�'�
�������E6�gOxVF<��H .9�� �*#��-4��}�	��� ��qc����޿��LQ��3c5Uf_��o���� ;���U{Cfh����?ӏ�?�����C������ ��'B�����/MO����&4�rq=÷�O�!�F�!���뎅��b�K��o<���ߧ����GT���{S�>���� �?��9Z�Oh�6\�2�q�/+K���e(�x���)��9m�m���څ����Q�<�� W����9��+�W��<֋�짏���?�ǯ~����u*�+蚍�l�H}^ٚާkb��L�d����c��u6U�9B�0�>h�ݚ�I����~;r�>���^ya��yQ�e��NT���Y��Ԓ$w�#��������׬�~ٴ��w�W�.��?t#��r3� �`��=c��=M��?*�TѺ�]��}s���FS�.�ؚ��%��7Ӻlփ�Y��[qO�a�>Y��һ�'dO|�-k3FG��V^@Y݁C�D}&sA��uu���3D��LՑaY��V�.;�	u�@�W�/r8�5�K���>��t�s��f{U��讹��N��ѵ-�z�m�fۻ}6�zR��tjЖN�	`&�5�������zMH�M����:�����"$O�%"<t,�2�� 6ՙ䊹J�9���;w�����ש���z�Є���+Qs#�-��7}�iF�wV(ig2X�J>@�Q������]����O���~�N��:[����gr���w�CG�l}3T�ti����k��ƛ.6L� @|{�%�5H�n��,&��uCQ�5	��ӟR�[�|3�ܣl��ʧ��{*�_�6Ss��g�K��v�+�Ԃ�����b��,D�LRG!a�~�=����]���c���w����{a����#�~����3� J���s���������Zmt^�jI�����~�G��vFft����[/on��9�GOt�{w��}+:惫�p�Z.ݞ�e���d"Κ��On�%�
�������ˮj�z��]ӻ�
�cI�j���ҿ==oU���'�A�G*��≢b���3Gy�?}��Ǽ��w{�/��/MtM��S�}�{{뮿��̏s���v�}�wc�����~��b���r޺v����Ll�i��[G�J��H�MCsl�eֵǳ"��t��M(V�rjVҠ���e��!�#��h�vC��>����!�n�b�
��kR�fY�k�&�%�e�v:奭���h"f�e�i�����~� a�C�_�N���|��M����н��wGbG/'W]�2�
�u1�$1c���&�ȾL��͙�7�ۆ��@�Eg�+G�P�YՀ8E%f2;X�G�[�j���m"օ�!,������q����� )�=H�z;�<����{��Oc�Mݴ�6q�l^����u�m��3c�QƄ�O3� �Μ�տ�C�	�1�f1������֓U�V��:�[N]�-6�X٥�n�ʁ�@"�dP
H�GG��mGL�&��}")�J�cZx}��V)*��ē��B��� (�=/�#�WI�߻-w�=��uް�-KF�x��>�~����Ff=��ޫ��Y�3���'H����՗)�^8J�5x_�fkۯ�O�t�Hf�K�����do%U�Q�"��(�x���y;c��P�����.�~��{TW� ��_V�E`�hL��|'�&������� x��$�V����{���;�ڽ�N�����N��z�����yLϪ��@�4q���
+Us_u�d��k�:��N<�9`5�|���%�K��H��� ��d��M�?E!�6�h�O�/�I���b�$T�c*y��GOʷ������{��������N��ٽ'R���5>�i��Ttv��n4��/�=��t�&�����ci:��hV+F���J
�p�i,��f�Qw]m��-,�c�]-C�sQo�򲙧�I��[A�$��J�-�6����n8zs��o-�PD�-dZ��[4�^ ���e���Y��U�`�0~�}���%������y��wmuލ�m���u]�;C՚�N�u���e\�--�1�,��}KJ�j'"����%c�V�֎�Yڻ^�cpS�^w�V�r����$/^V1~�H�N���H�x�H��] ٚ�F��Wvo]�m�t��[vk���M9���fb�Ik�n��9���!�Wq���|�%��ׯ�Olz'�-�1�������.���k=��zuom�1�a���z�^D�S�:GI�(#�Uj�ѵ"`��Y������hI���(�+=�B9����W��ù,6�֢f����mi<|!��s��{���K�s��k���'���δ��_�]��]?��Q�MB�mw���:�Q�k�]C\L֋BQcC��<�Y��h{����C���:��m���\�n�=9�ػ^���8z�,�#vP<p|%�)Q�.�m��~ꖩ��E}_L�Z�K���V�b�>O$�39���0�sy'H��}G��n��M�y}��7��O�u.��"YX�YК�n5�5�8�Jf&_���	�3�ᔏXo�7\zI�ΐk���o6��<T�;�Ig�8��(�QP]�,U$H��̻�]�O���k��؍tXR�3��ڒ$)=w�^#���c�}��m(A�5�e�Q�ߤ�^��@t�WS�]s>��������ꞧ��|��Y:+xYPN�����i�V09R�f0[$Eyc�v։��Y��:����۹#H�r��#nLB8�("���!���棫�^�d���QUc�]kT����p]�frY�{������;��5��WjI�3�4���L}6zoM�6VoSj�����}�{��hz�1+,�u�S��q�S�$ҵ*����H�#��*΄�V_�nbnP{n	<E�N��(I<�N
��n����e���������mk�]?���v+����|I�������3�:�c��]K�:�?��F�)�d`��k�;���!�s����t��g�,�(��Ôf�2Fދ��*��C0�]����؉L����@�ҩ<,�����*	\���������ܮ���Nh9}A��� M�s�=��K�>�ӏ1-�������pX��_5��Xů��,�����׈F�"�H�y'��������������$n�_�~���P~ ��9׾�{$���bX}g�A�?�o��?'3I쎝��_�wc5s)����P�N������d����Ij;O$ܨi6�^ɬ�I���{�� `��e-���#_<� �i�O�?��\�`�o�������~�0���}Q�=��g�z����]�c�fi��G�(�պs.��V	��4��?;�c�IweGm&�>��V,S��xa���n�A$�X��r՜*Ό9��O�+���a���9��y>�=�깽1��j]��jQ���q�w��b�K�蝋�f>���M��H�x��j���/Ùw�7�PU wJ�I�p|��Y���������2H��nU_�`H�A������wF
>���=�u'v���s��]�i؍7H�뤜�\��w:>��=���$O�Ԏ$)�����y�e��WZ�5�$�yy������=��Lj��B�O<�'�|W�dX�AK�P?ǂO,�~	'�����n����.AX��o�5�ʨ��{�9SXNT3y�i�Н�
(��Nd�~�/� �9� �U/��}����>N4�򅭓%k"s��[pU��VU��Ϗ-��Ȁ��s�.��&�$i��ll�5*�Zƕ[��*���LdG��Qه������1�8�P���2o���6�W�q��T*��I�tUy�L�ASu��6�U~�����Γ��8��M�q3UeU�l�o:�v���F�E,c�3P�&�po��T�v���b�J���/�A��E�Fb�� k�t[�k?��Wuf����qcf���4��$�8�8�-��%���
���n$zX^qcB�E��1�O�S,�;�`p�fZlUJ����M�Ҩ�\
�j�"\��[�6����\}�p�a�2�LA�i"�zy�Rm*��Nk�!���X��Z&E%y|E�EyݎY�Q:Sb��8l�Ԩ*D�>���U�T�2��P�9M�������Ȱ_����=1�3fYJrM�pF�E��\�a;ۑ����]�[�C�ӎH�����T�V���*iAB���>��Ɣ�c���/,h�8�1�VVW�hYx��߉���<vf2�.�ny��檳���6��K�� �ʠA�6c&h�j=�� h�-H��$k_�f�AR1}�R�+�Vƌ��I���%�&�G5������ �P���p��+�?�$y
��"%�P��`��cy�o�ۡ�G�ё����J�J! KƊ��Uf��T:��U~/ͨ9:��t��ۋX�"���S�_�y��E�M�C��g@�� ��ce
X�.><��;�2z#5S!��,�Yn�����Fbfc���NO<�'(�h����oᒳ:ő�`x�錢�21�f꤁��k�*�V�3j��e!O��em���99�	���u�Di��!�Z����:���7ۈT,a�Cc c�|�'�]jMR��
ұ,�;����Te~G�Vh�/X�c,eDr�<tly�CSr�	`C!�U���[��^3ΠFi7i�^j�w%�F܃����59��!�)�AF�p^&�p�_�ԗ �P�1��88��*yc�nǑ`	;� $��Lf9����(+��+^v�c"t�6u$���ı�k�q�|`ov5��4G��ѩ`X��K>�X����<0��5e�D������72 �#�,���ub��˺�cZ�����vŔ�h��gd�c0��'ط�N���n�`%b�)�GQ,�R{�_ɇժʊ<��~��Ǧ0P4�`�l���j�;UU9ͦ
�W��+�SGp���Ui%����Q�Svv���!��x���ʇ��JE�2Ehݕ��v{S�J>6��5x�ۂ�d�켋6��EjQ�M<Ve
�0i͟��m��c����U�R�1<7(�^����"��-T�~b���C*�b6GT�^K��o�U��z�b��jW�Wvb�܆24���yC1Ỉ��$]�Y�<��-ُ��r�U�� �c9ex��n�+kc�;��F�9�	Y�z�!*`LiZ�z4���(�S��$��^c�v��5KR���F�ѧ�� 
<Rl���4��vv*�1|jG���h�+,H6��=8K���Ryq$�UƎQz0�	㐐�34f�L���vg
8���*���� @꿌�:�J��"ě�X�.�D���+3V�`�� Ynܾ9�,f�w��~~)8XЯ�tT�#�aͲ��3�E3���3�Υ���3�����#��m*��c�����+;�-;�3�-���ӈ-/6�=1���/o���گ��P�g�ʅe�*�����HnJ8�x�*�}1�O�_���1�Ν�5.��.yZ~��d���:}��F5��R�	�� WV�F��ӵ-CG�_S�oK��5tS�#E*��u �G�_j��=e��i��Z^�FKM��&�<k,2��̑�*��9��H �;����}�8]��c�ש�C&������i�i�DH�'�ty���3`K�:Λ1v��ԛ{y�ߐW���M_�B&�`S�G���x��	[��+��Z�;�ȻE�ze=�"'ֶՙI4y�&�N����nw*����_���q~�s�=7����T������zo3H����4��l���ᘚG�}#%3t�/)S#/v�)�NN��b6����v��4IN��u�'�f���O��/�k��"X�U�?c��5�~h�������^����<���A=yU��d�XTg��{�rwC'iv���v��>�t֍�_����Z��h}��ݓ���=!�dcdOF�N���S�2'<6�:M\�B��5Cw�l� ��Or�ߨ� �wF���~��)�,�;��Zj�"kK4rB�g�ex]e�S����-���ُͣ�[k�_W����F���HR�y�չ�X���ճ�Ȭ��t�Y�{���C���#ۭS�ݑκw#�������T��Et|S���i�o<f���tT0�B���.8ȱٽ����G�A�������i�X:f�Q�Bڍ��i��nʠU����!�
�� �u�s_7wĆ����lt�`鯢��j��=N�R��5l�Ez�k<���Z��<�Ɋ6�Q�����=5�oH�f���P�v��Sn��Z��霮�ֺ�I �<��j��k�/c�F��Z�a�"���i_�i�cp��t�E��t�pK`!n��S]�P���ૢ�s4��9�i�~֧sUע��-���HC/���Jb��Adt>��ܯtP�ѧO؟������{�0;_�����ް��gO�����g�po�c��;��L��0[z���ۣ�qi]j۷��ڎ���y���<�_��^h�d�"Yf�Af����
�͑���������k�:�Q�]*�.�r���Oei)	b�0��∺Ab��eιw{��W���]��{%��� �ݯ�zB�]�]���{��^��Ğ�����t����Z~4�Q{]#)�ZIV���� L~d����$�4�=g��B�6�H{Ng�#ٵ�x������won1�� ���򶡶6�س��^-I�ݖ���KEN���M�BP:�Iߏ�	�#����ԃ�=��Gz:b�pLmsC����:�E��m�;q��=A�gQ����y?hN�8�7�U~��	v���z^�T�*ݖ\�'#�k܆�H�����/�쾎�� k܃q�M�{nj�rVh�U�Wώx,LE�[��0H������wO�.���0�ߵ�p}���e�̞�u�oNv˻���ӳ[�r��5o���r���|�S�JҬstu�s��3k��Hz���Syh��OO5��Ӧi�	a���&�t�:�õ��X�eA瀼R�<�GG�ͫ�H�]J�2��P�d�M���v��a�}!�i�#�DI,�i���A|�;����]]���"t����/��W��^v����&Nv6_���Ŗ6�QY��n?�Q5M3T�CO�V��b�KH��bH#���o|r��1�����R��n�bk+�	�����Q��,��=�F�9�F`G�9�:ο��ε��Ю��XAt�.]G��3��4Ҵ�4:cR]UV�Zō8��o�6'��ёk�^K
{��~�=�v�����pO�25���1�	b8�"TnQ��
��>�? ��{q�Q�~�{��}��t�Pw�u�Z�_B�Z�Vgt�HegNZ�[w���z.�U�2M�V^*O��t��VƿSǣQ��Cji�1R�h㑒�C���*�kq"��l��־NH��MVK��1����tV~;�5Xcf�I&��@y�Fw��}��_�W�����^�t�}m�i���zh�׵��i���Fi��ֵ��S��b�j�}CN�l9�pth֔�z˻SgRꦙ�m�z�l]�1�A�D�\�Z~l'��fWU%�R��Kd�"�ۺ-쩴�ɧ�o=���5+?�.&Y{L���uT1��mG0�h�HH�_���=���^����{��*��}��fNuV���ftOz;��X8:n��>��gŢ�bK��X�"�����tx�k�����t�ըϴ�)^2ٛ�4������/��ܷ����D���E��.��}��7o�}6�-ů�Z�d�+�ֈ�Lg�1����N;��~U��m�tG�=�^� w�����/|�_д���tl�tw�N�ӽ�v�AǾ/G�'TwG�2)>�k��Q���~�.�Li�Bb�mк�Э_�s���i=I�rI,j�6�S�If�az����li՜v�Y�R�#4�<-U��u�]	tk[WG�:x��1���V� ��dԵ��d�37�fz%�8TC�T=��I��_��G�[�� �)�݁�������v�'\�Κ��M0N����;n:�@jE�m0�eFy�5��"��Pl7���N�Z�{󨚎��k�.��K��
���e�L�&���nB���6�p��B�fސ�Im�lz;z���w��$5-EZ�1�Zo�W4���򬱴uё�Qh����$I+��n�Һ���o��������?�]Cn���z�Ϧt� GI��,����5�Ϛ�V�r4�g#"� Cx8�ԭ������>u����kW��7H�[֯�D��\�*��x�G��ye9��b���>&�C�ޙ��ےX�[7�.��l�v�ҥZ�I'�,���!��C��v/F�&����}� {G�#ҽWTǿ�n�'���]�u�`vˮqz���l��=LfO�Z��Ȑ�􌝇�sy|e��}�_��f�����Ӏ5��'Xӓ\D� }F>`�b
���<�Jw���-��Ս��K"����4�GG�>�d����KNR_�5
�`c!G��P ɝ���폽�� �ݫ�w;��/l:~�zk�� Ow�4Oq}��I���t6�\M�wC�\'��|'��5ӱ����'�A}L�|n�kU��� M��o�<���Bi�9�4�,��^5�ևrI���jL����K��c����5=�.�;dM���STy뾏zD���R(g"�2W�!��,D҄������K�t.���n�w�@�:�36]C�>��&���]�]3	GQ���;M8��mI�)�ӱ��XqLvȭ"G��Z�nѴ~����~�
����GJ{"�&�VC$z�����F�����Q�������w���˽�O}$������$�`�*�SP�%N�=�eR9��bo;پ��>}�w��ݶ���a֝�����z[�������2�ڕ�=}���awp-?+T�Ǣ4�Q·"��㚗PaҶ������1�,ߧ��|�5*Q|�2K��q;U��y�@y�~	��b��ں���%�2�\ѕ>ZPdX'���P��X�̦6�U�Cߛ�ݮ���a��^�v�����)��n��w�z���i����+�_U���,�Ի9�d�Օ:SXjc��Q�.���O��xn^�i:D}YԎ��i�djz��k��J��QE'���E�B*�����%��c,`���K��Oh��6Ʊ�D�4�1�����y�v��M�X7��dI�$�>N���mtRw�]��J� o~�:��һ��C�yկU��sz������k;T�V�_��thxك0)L|��q�1�op��N��3��*�Z���?Ul���*5"�Ql��,�X�ix��XXL"��g��l�Uw���M���O����ӏ��5��?l5�$�멒PD~d��zo�5��ܭ{�=y��Ӭ�ߠz�/�:���^�,N�n��T�V�H���������,|�z�dʮ$����`� �5��=f�T5�(E3D-&��Й<�Hl�I":4�Q�蝠؝3�<�����M�h� ���):5�FH�1eY���tH!�Ь���Gj��3m��u:~����^�k�����p�3n�tg��t�z����]r��>�� '�ũM:�dC'����!�B�]�l.��6�����u�mS��;Vh+X���M���yjH ���� Ǩ��R�GQ�ߺ5��osip��p>��n�be��-xlD��`�����H�s!z�v#���t� H�m�{ܟu�#������K�on����;�Gb{}����]7��Z������!���P�q�<\�>���
M1��N��:�͟�uCmi�o:/ׂs0���|^j�B�	���0���,#V �+Y���� Ww.����N-�Wu��@i��iʿ���gS�w�vA3��Fz�w{���<���u��n��}_K��� �]q�mw���]w'E���~��l�m���qRZ�5��V�)c(�Z�<�O��TuMѬi�]��	�V�i���H$1O
U�7iQJ��r^��*���Cd|t�M��j��Ж[��47���w�K`?�);���X� r�)�j��u֑�u�����.��^��绞�=W�����������.���ݮ�jsl}n-����[���8�����M��n�E��SA��z��f�ӃZg���]Op�<=�R��BU({+_4��ס֏�:~]�opصZ�UXM^W�"+1�:�S/�����'�����s������E�K�=��>�����?t{��<n��ozˠ�K[Y��>j��rƘO��.6T2�a����a\�P�_�d�Ɖ���� ����/b�O�yjG�V8Qʸ����9�#�a�6���+	���2� S�q�RҼOY�@��K/`G�ɅY��F#'4���Wi�)�����z{�=��ޘ����Ǿ��9xz�Ui]+]n:���u>��[fc5�^�lgԪʘ8=;��_Z���V��j����7�g�j0���򑴋+5+h��*��7�v����;Cfĺn��54�,^Q�s)ɞ�V�FnA%�Ԑ`l7�}��G�n��N��X`���qg�����F���g�n���Ε�Z�MGM�D,�m,�A�K�z��Ae}:d�J@�ZZ�G�;�A+�YpA>2�Ve��V��E���ERG�����&9Qx�o� �Y�-w��q�[T��=�j�G{���3.����Q�{{�ؘ�x��.���y֦v�m�ΏJiT�ܨ�S9t�n������3ؙ�i=�v�to@�"�`(����Ϲ)�$�(�$)�J��>�I�<���q��;�g�a��t�����ߑ��W73R�A�?�]=�!���S�?@�6?����tl���RNfS��J�ؘ4Q�J�	*	%�y@����� <��x@;G'�����=��gT=�{N�'���twt�g��[�תu�o�����iS�I�F��j6��2%f��������"���j�"Kd�V�u�Z1����ڸ�=��cvR@x�n�
I=��Kp*�	��8nH� �n�
�����9�s�ݻ��l��vL��}OɁ��2�s���R�#�gj=G�eu	��m����8P����*3�ޭ�Z�?{򁒳��U�F���$�z�MǧQ�>K�W�<f��v-��H%e��ǲ#�����gڼ}W���v�7]掳���ڞ�����;�z7T���o��>�|ZKJ�K���t�i���&�JCE�����cP~�$�$����/�R&���Y���1ol�z�v�2�����N�{��a3���6]��S��?��bv���6�F��6n���#X�i��f�Mr���	�%�'����?�� ����f@`D�*�1w��>����5�d�Ŋ�ݏd܀C}ى`ă���a�թ��H��>� �gǙcH��������$*�9�F� +�ܟ���|�	�p}z�&���O����𮲒�뻟�˕�Mu�\MR��U��Pg�� P�R՛m��� ���a��j"�!�����O����B0dŘ��Q���� ����B�5\�Jzv����E#��x�E�<b��m���?;UiN����H��������~��sY�O% Y#?n~��˺'F�A���&���ȶ<pT�kdyʒr*Y �, ��o�� ףi���l+������� ��������^��������<={�G-ZƷ�ɪ	�S^}G�%�q�N$�2�I �UEt�p*8�R�c�5�,���9��o�����Yu�GҾ��y&n9=�/���� _�s���n'E���5}Q�;�e;L�9s���TǍL��Z��+�6>Z��譓2������uN��iϦ:���~�y��P�NJ�2�b8��r��J�+\���$Vf`܅�~	�_QV^�X�}+�o^�:'�4�s�����~�{К�Iu�_���ھ���i�䦧�+�'��_F��e�� �;�m�L�S���G�ɐ��6gbt��;;]���mǢ�ڋ�i�3ɧ���T��*�u�J�R^
H�!�}�ͤ\]�r̶i��MI+�x�>X�����l���F����������}�� �"��.����-��G�_����z�ii~��]3��[i�3�t�9f ^B���:�砛���E��j�R��ӭ+iݳ^��SR4��X�0g�TkZ��Ù|��Fd(�>�ͮ��*������B����^'���lH�G7r@����R|Q�2�2�\7;�Σ�6��� ۯ��n>��~��;��#Ӗ�>u���z��d�_��.�E����;�M]G#]���ɥ�u�l�P���@������fu�\���:F�5��E����S�x��rȍ��4m4��ӽ����iv		u�i��tw/M�.��uB$�k$�KU#�1��V�j��3[�%yo4��9���=��/��W�4��s�G�_py�=����w�]-�=���չX>ms�;�����Ҳ}�j�V��h�^H�l�wm�����⿧l=b투0��R��-sZ���Sҫi즒�G�If��A��;�@�ת�޵{����k�A�i����4�Ly�1>}ⓕ���/
Vy�3;��ﷸ���`����O`zgއT��������G�{~���n�̎��;eѽ�Ҹ�Bh�s��<}+MN�gy�|����~쎣k�2�v���ޱV�^-ǧċ3�Y%�wSbku�-K��y^ǘ��*�]�����hP�W�h�f�J��L�GjiZ.�H$��j��x��<i@Y	%�Z���:y�M���CۯJ�C�W��K@�� z{��^�u�w�Z���.��j?��ײ#sAl��7���ϴ=J궵�k�^mWc�^]F��ٻB�������
�2�v�7�)@�P�>16/K�6��[�~������fKe�$��E�����W1Չ���_�.����v����zQe�Н]���k��YZCL���SR8���k�&�O1�pP�4h0����}��iz��ZXiЎx�߼�E�G?�U�O� {�n�S�z�ykܹ��Z]��I{�=y@<v�]�H�r9*�wE��؅Ϧ��W���t�n��=ѽ-^������{A�l�� i���Ѡ����u~N=q���Ul�7�Þ��Pm=����[����sT�cQ��؝�Y�?�����5���k�3�Z9�����\����z5�l���v�z�f��~�^� ��狉��@9H޻��r�������/{��ߩ6D�G��j�L�����=��}M�b�x�{�:[d�:�fs�';
�͋�$�/Y?�˖|��k��mG�i�,�~�����Ld�u���N��ՙ)̝� ���r��G�[�i�1��
}�'Rw>��L�ܪ؎E��������w��'C�X���w�UUn8O�wGX���)5
�ѵ,� ˧k,N�#A�t��Y�h��Pu"}�6v����6�������\���?o`�?S�7G�l�'9�O����-m���0�َ�������ɬH#�_%f�|�`)�k���c���_b_���c۝S'3�?j���t.��K��aբ�M�=_�Ʋ�����R��=�b�|�\G�F�����=_�wm�߲mM�m]n�0ݦùi#ӆY{c�b��O=ILHMpHn�|n^���Kfo�1雗B��b���m���ׁJ��,��f!b4#��J���N�w����]����'�]�w��'���ףt~�h�e�-'ZM.��Fd:��Q2Nj���ɍ�'2���B�g���h�V�=`ַ��%�2�ըݬ�X�\G����e@kH��d�'g�By+��ے�N�{c[M6�5%���H���G%���ޅvo��Hddv�,qE� ��<ѽ�{����[Ծ�;����v2��w���#L���Z:�p;=��a>��bY�Ι��Ϡ��#N��=K�֞��Jm?N�==F�-��l��2W�V���J���ֹ$�/�-U̍3��T�ZtZ��ӫ$�K-��z�eW �b���M��>Xa�c�wKRs����G_�������]�8��n���ճ�Uize�ǢC?[�p�m/�]��㛮.n��j;`[t�q�^U����CF�RugA�w$ۖc��o$2*�XE&���w�D߿v����2egf�W�F��t�aT�u��R-v��D"uI���]x[��d�U���U��H
�(�K���]��Mۗ�/���j�SѽM��j}��:�P��h�t�S�h�ϧS�=g�0˾��.,��(8��M3KHa�:V�"h�Gf`Uc!#�O��Xdp����pF�ٖTy.;�*;A��GҀ�yz�p��t�ۯ�<>��|}#^��O��Rf_*����������=����ӱpG�$?-�K&g�dի��[�BѼ	dX���B���q��}���*�)���,�6���>3(������q�pc�<�P'���G}������>��/������z[�:�P�4�l��������z?�v�N��V��I��5�T7N��3/�AR�5d%�
yEy��o?�Ǿ����eR�5�2�� �^א��F� ��/c5�״.� ���Χ�:n����h�� �;������O��29��~��:�e'�z���Zzv#djyu��ʿ�M,򈢍�O!�}�Y�����>��>B"/,�4���?�����}��M�Y��n�ӻ�����Q�=���=5z߹R�<\��-O��)�Ռ�s��]g
��
�m�R��񴺄��p�v7�� �9<�O�I�߮,v���Q{���$��-�<�#�9� �l�W�����U}?U~�w�S�������iq�<���]:��M>95VO�9�� ��,i�h��m-�����!缡�I�)��O���?����j��������) �����P8a��������KvGT�I�������G��ZCO�Nv��]'�f���}5���Һ��z����}��Rm=��6�ײ�d�L��ye'�]�����lr���$�_^H���d��ز쪗E���J���>�P/ܣ[����=��G+���ެ�>�������������z6������FhQX�;��;�L:{G��Dd��H�M���Cj�ʻ�2��}�'�<�I'�LĳI��UTU`�� �z ����  >�f�f��t.*�9+:d;y]7M�6Gm���$����G��qA:������r �?�n�����~��~߯�s�C�昺�Oo������ɂ��=���][:�"�sprG���S2������`ݝ���@����?bp෾IoD}����ͤ����Dw�5��v�a8�)4�R�6��<���74��2���%�W"���������T㎌�2,U��Ya)+VB��Lu#&�|Y4	�Fa�f��~N1ݸ�qc�+B8yh���� a9��	^n���3��]�U���m¬����d����=	mԲ�cɌ��?ȝ#9��i,���T��*;/��P7
���*�V0L�iUEQF~*�Ũ�-�G&���W�Q����V��.\2�%>Y��� TM��B��|���X� �eP�6`���r���1��`�sD��ȅ$�Ɍ1g-��{�������!��x� ��O�'edLDM��q�J��w��ob�HP*�[d(v��i��d ��Y�Tx�d��r9���T�y���-E,ܸ�7(`ı�,��w���u'Ɵ�4�d�jJk�~Su �=1�>r��d��n�2BP�����&o�K'�����ޘô��x�Lu35&y4R�$I�"�C���UP��AŌ<���F[�=�gqN4f(UYZ.�P.��yrm׎����&�R�U�c����ǢGu�%���T8PWv�сc�\�hF�J'���i��9�� @�	�U?g��j��:m�`��YL��y�^6E_��H�ITĳ��Ny���掱�9�X��KyM��������*#���_��3/�����-P�o�W�X0ݘġs���m�kƁ펑�~+@�+�� ;�۱���q̣�]����2O��փa��dI���I�V1�Ɍ����S �ɓAi�����b�[���X�_La$)�Q�ŚBE]Qr���$*���`?W%+��,bO��o�0F�^s��UK@6����	�IUyr.����ʱ�I�}^����E�"'�XM��u5p���L`��R�f����9�� ػ�o�l��ȧLed��Lu^s2_�-TCl��j�Ѿ���K��J�
kU��`E(��8��Hд(P8����_rA��G˛^֣e%D��3$�+TQ�l�-M�>��v�1�l� �B�?�'`/��L�m�G���Ɣ�hV��1�3Pe� gi�U?�KruU�rN^�s$3Dwa�%!-#>b�F�fٶ(AV;�����>[%c�$�)��Ndϑ��f<S�����%��B��99m@t�������/�3N;�٬�q�e�� ��ɤ�������g�Y��g������R����Ō6F0���K�G� ���Eevy�-@~��o�"���P՗��j�fƭ���h���H�W��ݐ�*r`X�*�dc�FnPP=�6|T<Qa'-]�@�m�g5��%�8ܲ%7�Z-B��!'C�&�	�Y��b�쌄��䱐��1Rћ�6�k� ���ނx�w\R�ڜT�!yrB),d�y.B�գ_'�:���$E&N̞B����?$1�]��A7U,��F�wA�
��!a��
@$�"���cM�b���B�Bdc�6��C �)��r��0�L�c.Y���2[��}������2��Q�ܱ�9�2��j)�*�O"l�e�ׂ�+V��s(� ��m�ʼ��ȯ7l�_+2���M!k�$,΄3�t!����9�U�Ym�@�V���gae^7f�ʼ���/�'v1�ʜf�X��fJ	�������-O �eb�7KL�2�Z�BR�t��'e`<վ��
��g�R�X��ÝOی�g��r`�� �ᨔ�0��e�"37ؒ۱���o��#]]HW*�ˉ�b�])���ĩX��2��U�Z�+-<m/�������}[A���}??������i�����WʚX�}��e�����+��O�����e��U� t |\T��"x��CA��lO��q����XU�caٲ3�_Z�3:[Sr�(Fv�e�7ǖB4-����9�]A�;B;i�/�7�YӬ�z�y,�X=i�"�f�N�ȼ����M6��jW�*�Gqi'���W�=B� @++,�Hz��j�n}e�_�b}�{��>�������bi��Z&��(i��T$�\��xrԦ�b���*�}���)Rյ�5M��x�%�H�e�-B&�+���
�P�/Z�}���on�[:WP�SsD142�4�3i�E���-6�+�-�����
:��U-��:��}�^��<>��龾�][@�N�ͮ6A���,K��1�/÷��VJ;����ߣu3h��.�әtٞE�R�|�Uya���j�d���גHgN��G,�+*��zM��Ce�Y:��=R��~X��M�1��+3�d-{Ѭ�F�MSװX��W�������{���|���d��n�hy��Dh]��V��vϤu}+*��n��ύ|��Þ�U���nS�S*I<p�J?�l՛L�R+jz�'�pl\���X�*Ǿ4b#��Q�b]�q�z��&���Z���=9Դ��U咝X�2q��j����d��	G#�	�gk�s?QOy�2uv���֝��&�Ӎ\x�tΖ�(�����!Kt�3Aơ�;���XҬ޺���g���7aҡ�}di���{5��y�V -��;P0U�ޥ��7_z��_�%����oQ��H�iC$�կjı��G��1�VVv=�N}���a�k�?�/l;5��h��{ܽ7>�:橇��[�h���u�w7R�1������r�����4�D���=8'�O�]����V�ƹ�.B��X��L���;�]#���������-5��U~��C��SmmfS�6��$H&�5V���y�������H�?"Eh��}��T{��y����w[U��[C��������zOK����si�������ޟ�h���ֺ�'N��3F��E^5�t�㹯j�㯪U�FRD5cht%I�t	�D �ߛ�X��
$�gi�Z^�RKz�zĝ��iD��x�>猕Q���x���9ѝ:���v�ܯ��u=��5�.��zS���1����Z6�����Fej��?՚{ꘫ�L:q�^2�]e��<u�n�ݠn�y,.�qV��3�={ �Vp���s�F�6F���`[nk��H�LM/w	�4}�Hg@�' �>�����GXvE{�쓹7K���GFu�r�O��s�x�.��W`��z&���u����z����9�Zk�'B������k>�k��kٻg�:tGj��ǤԹ_R�-�[��k�NZ�~d
��_0�,B�6s����zi�u�'��3K�,W�VR�R��s�O?�v
���TZ'R���3�^�Kn�h��{I���k���U�k���oW鎯��~��M���L�����p:�SǦ���������328��	��u��� W�66���Z���(��3�*rͫ��4ď���Vy��F�F��uJ�v�}nr-�U�&����Ga/�V@#�Ii<^et�	3*�RD2f���{ǥ���1{�v'�Z�r��I�0+��i��\�'�^�_*�zFx둑�����/��v^D�m&��M���U�]W���Z֝�H�"�V��uWD�UY�ǅ��s\� ������}�4�odS����y��ࣗ�R��"WE<�*b�V6n�c�˻3�'��n:�>�s�s���r��G���t��P�����SR��c����^	�ݎ��`�c�:��:2LP���'����� X�7���i�S�lA��":m&��bwGTmB�1��ww��Y&��)���9!tצ�IZv�Ι��Y���amF̈́���"2w-z�K��BQ�u� 2GM��#v+�����Qw��u^��{{��d�gPtp;��ך.F�t��iY�;Ӭd�����ʮA����K��ٱQ_[��B�X�9���]Ѷ��
��ЗO�(Uޜ�sh�<��>=r�M�u��%f}�~�L��S{�'AcX�u�J�+c��j��.�4mT�WN��VMP1���V��W9�ێ�{f�w�����O�~��S��S鎚�����b���y�;�`M��&�g�q�ci��G�&���n�ڇ�Z�{؟}t֣�4��]%�/�:�M�b���h%�yl��H�P�FBClF� ���V�Z�ў����_p�k]�lWH�i��ו�X�q�ahL=��OE{��W���$��{j��ҽ��z���:�Y�����R��t�68�Gl�
��;�'�`4�S��# b�r�c����S�ft��[�� nMoB+�U�!��$��:�ۑ"�d<�HEB�*#,2*�$}L���:����L���^��Ȳ��KMGᆵf�ު���*��� ��'1fY�n���O��ϭ�������3/�]����V��[�]]��5�r�r?������G�Q������d֡��(g��}r�_v]���]GV�t�c�i�>�43�ڼ3G/�R	L�e�,��m���F���17�;oj��t���+S��i�%K��
�V�5kr@Q��, Ԑق	V���$o��R rc�>�?M�a]��^��^����C����}��o[�{%���T�mP�����N��,�������<LxO/�ex{����w�s��:���OK�5�`�-Z��DAl�� -#�s�Ě@H���:���>��"������ ZG0�5���M԰��宭�ӇR>��pD �����c�T� �{��+���{u���1��=��k�Ȧ��N��\~���r㘶L|�&Z�r�x[>�����w't�@���m��n�Ҏ�������~T���m~��r"�e�H{ǒ�0�k�����Hڝ�7ņ�7S5B���N�H��:dC�#�Y+��	�Բye��X�H�"z��-_�#FOx����v�����������ף}�tD�Zm0�4�� v�+��钥,�+�1��L�'';*-�_t���~�Ao�[R�{>���4]"=I������ �$�������bb�T���uXOnN�M�GG������w��:��~z���k��6W��W^�%̰Ze���,S=���7��{톻���O��{��S��wH�'k=��C�O/�Z�d�-KX�������H�ϩ0�V��G	�I�,�=X�u�A�����گP�l��H��W�ǁ�%;�w���D`�[��B(ˮ�����~���ې�ݨ��:U�M��P��6���C5n��~��/w�#�y{��7n��w�T���鎩�4^��~�h:f��ݾ�<g�(�K���/H�l�[�Kc5��l���H�ffd��Z�/���m[��Z�<�&�P۬�$�m���3�J�9$e�8���Q�ie�:S��/4]#^��Oa^�[2��� �w�xF2C����iIi{���ޟڧr}�wK����폻����Դ�u�@��4��v�K\]_��G�\�ؘ����|O�y��t��t�C�Ǵ~��Y�oN�'�m����gK�=H���S	�t�$xm��q/�W�Y��4rI*��T�M��Z}$�ƯGG���j�6��q�UuӮ�-�>b�Īū�6�b��a���+�]�������7�y]Q���zǪu���;�ۭsM�z�v;!+[�s1O"���l�X�b�%O���h[�ju^��<��+,7�?>��L��^^h�A<��ܫ�������O�>���D��v��⶟[:<�����E���Y��*iX
�aVPNj�V��r=���;�@Ꞹ�.�N����j��u~��q�B4�M3S��Zh�U���Y�ٸ�_7.Ԧ<���i�:].�t�N�Mx�=�A����mזx�B����g���bX�E^.�{�^�tU���'�=E�K�-j�=3�ZT�U�*�*�Z�3ٓ��H�<��@�2߳~��<=���r{y����s;���7�����Ժ�D���ղq���.������Z�uLj~"�!�#S��1l����ϩ�6�Q�"�iܥP��GF�tH.���*[�6�0�'��|l�����ң�H~N�W�]B��*��Hd(|�0�?s(S�����{�4j]��i�!�]�=�����{��E����-��g��]��c\u���=1~+�y�N[���tP���[�h>߱0I"� �i4�����ܭ=�9�'�m�b�� ���K��Ru�I�,m���c֦�W��l�anK�X3��<55/J|y� �=x�f:u�w:]0���{��5.� ���*��g���r�O��rU��K��Id�j�q�y�D��>�Ԝ�cG[���fΒ�L��@���5j��[�o���;҆��1�MF% )
r���鮯�柨={��ڷgn���aZu�K��R/#�# �؟�C�+p���~������ퟬ:+��S�Q�J�Ƴ��%�zƯ���ع�?��|l총n$���n���11r?o���2^կ˭O�[�5	f��$�;ܑ���W�y�?�_��� �تB��V
5�W�4�1E-XՔ8T G���jr=HG�ͮ��)��gp5���A���Ʈ�=y�]K��L�Ǧ�+ck���V�v�.��4�\ɳr�<Q�ӡ�Q-�ܺ���𺰫"���iTc��C�`[ь�� W�.ON��r�O2�;A�'�|O��`=����wc޷Hvo�5.��7l�˶�}���u�4���g�gk:o�^��V]`�j��_�&FE� .@ѿ.H?V-ٔ��|J �T��y���������p�"p����]Ò�� /^�����r�J�#�uN���˗�i��F���R�9z�-s������ɦ6nL��ٍ,����R��Z�'I'��I#�Q��r�e�����/z��Փ��X��T��@`O���o��ٯr=��{;�Q���a��.>���sR}7���5��X�:���>Vi����E�\�^Uq��Ϣ��WEI��=�����,�%�_�BCB}�2(�<�2�+:�a�mMKr������U����)x�r=஗����`{Q���NӤ�Q���I��Κ�^��+H����M�;�����,��Ȣҹw�,�\Ɯ�{i�����֓Ow� ����ꬣ���h�6YY8���<�74)��IdG�UI�f{An�"24�v9���g��|��-3/���z��z���>oz���� E�V��J���vW��J5��Fj�u��).��L�?H���zMWT���������ݠ�/�R�'�O'*�i������v%�eB����K��M��ƥ�Z����O���I��y�z���k��f���ڦk���u�[>���5
?�ڴ��@��Ԫ�`W�sq� ����go�q�
�����N�y9x��z+:R�I�u��~�f?�� ��c��(Os'����� |�{�`���_����:$s]^��.(�8�J���[�������w?>�$�#�5�bN��}�?��U�G������7ŋ䍧�d�%�o������s��($�w�꺄7@И�������Uh�$G�� �{-�5��beG�N�V�Y<���*�n�6��w]���	�G�6���G��|~r����T*x���>�-*h6��g���CK���xrg��Մ	��_����V�GU�A�:��K���C���>�#��}����ek\�QeG>��{�{�s�������ִ�����30��ײ��i� M����4��Ky��0; � ��F���P��>�B4��cd��Xq�!�=���� w�=�nҝ�jY�	�;�����Gc��Ǳ�ْ}�v�D�	׺� Ci]���e������4���;O׺��3�?��0l^���b�R֤�nu�q����bӖ����(��n��-%��i=D�u�=�,(����-1�#}c�#@��%��F������h�@i�C���RJ�0~�`s��ʽ���p��ܧ�_�;�=�������}H�KD����/D�u�q����{�VŌ;9�z�����֎=u���M�V��q�>�t�i�΍T��oY�d�<枟)��ؗU�do$��h1U��")V���4�'N�z��lh;�Ui4y��e#qVt��בx��iD�&�TX�E�"w�?t�{���ݏ��싨��뺦NL�{����oq:/������u������&&�i�W��E��\��Һ�O�7�%%���M���Re��Wү�7c$�#�%����X�$V�a5΄��Ғ�m��Q�$��z���*,U��2H����I �Onu��z��:޵z�r3}�t���#���S�{T=��S��fei}���^��Nһ񕏩(�=��7�j�W�� �A]���ޖ������N(om�u!�m�?&�P1x��v�JE��r�L��V�(�PG1�$j|;�}hZ��ڃzZ�4�3ƻ��H�$�_P�b9*[��"�,�Eiͅ>HOpv���ޏo=�{������j]����u���su-7C��\�+'���'�b�K�<��B�N&��a�ul�	��u����BzE>�Ҷ�3R��Ѧ��W�i��)KdO�:��ΑԊ�֚�i�,���ˏt�:oSz�OlY֬��ڭ���)�����P���
�7��U�y��Q"��v�ݷpz���O{J�ѳ�W��W�����;'�8�{ۮ�n�����'P��v��O�c�&fvVvO��M�/��gV�������-��[���ƅ�X�>n)\!�j�H��#덡�k UT����~鮝��4�t����t֥8@J�X��O)</cI/,��bxӿy}Q��o�^�vK�_�n��÷����K��]�O��s]��s�~��t��?Sdi������c1<z�޲e���z�o�&��d��v���,C�V�C�<0O$qZ^QZ%��3���;��2�:�5ޔ�\Һ[�O��a�J0۲����IY^','`#�	�8�c`���%���\�����&��������:�Qc�'SwG��^���Tw���~��Ե��-�e�F���u����žV����euٽ!ܵ:=��ۺ�-[�N�:֒�����H�W�Z�y<Q4�+/i#åz�����j�Rg���dʰ~�yf�_1wU�v��"���зk�!B�)�>g�/�cF�7�`�!�C������Y���ڬ!�����(i�]A���8�5�:mi����EAC賺�7�i]Aꕝ�$z���X2�xZ�唗��E����$���G1Hxu㒫�9��H"��KOt7r��8��/��F��r���`HC(� �e��R� S^���{����ؽ_�!ӵ�o�}K�t�s:�E�RѺW_���z�E�0��V���?�-Jh�ڎ�T�5~�G��+U₥�֪��E=+�
Fc��V=��O$q]���T@�|�:u��zwU+��z\׵�b{�Jy`�VؚUu�b�<�@"y�J$Dv�<� ���y�����oݖ�֝������ڿY�[C��f�m#=:���]kK�t���l&�w�?�^������ͷ��WV�n��=5ZZ>�
��iS�d��?�M:�^Ěy*�8�Eps�+��v���u/jA�jR�����+�Y*Ha�V{��2�;F6iCKX$20�վ�'뉓���K�-W�u�o:�RjG�����k�����~���蚖FF.���+&�ɻi[��u�%�z�or��*^Բ�^������W�D�X�9q KQ��3v�}"�Bu���VI媒O*��-�9��x0ՙS���������� �WZ�{;_�>�ѽ�u�.��o�J���u��JG[�}_��u��	i�����rU\�<�hgQ
��4T����Y׷��*���.ؑ`2�����4�x!�<����?�	F���D�zH�Z�װu���@a*����#�mc�I������i���d}�u�`}��~��t�'�L~�h}�������t�>7_h�HdS�>vH����+6��t���ڢ�]CD�F��������{�ڛ�M�X��؊��6Iz�/�P֩�:���D����&��~��z��7��}t�:�y�Ժa>��2��!�����k �f����w���������tN�b�ct�Su6���v���X�~=z3��S�2k�u?^��o���Q/�����uEƟ*4]b��GY�f͂D4��U`�� ����#�Y9�ٽ�z���&��ҡ�ק5��N�3O�s$ӿ,����|,h ;�������)�_Ku��ju�y��7�Y=}�n����i0Ӱ�ѫ҉����x�����š��u�f��V� ����]�$
��d�C:��I���e�{�##KVd��4߽O!'��cr� �*�����~}��~����C�>�t.����GP���]�v�P�r:w:�Q�ģ�n�<����zfưz���-��e��&�槢ҭ��ӵ�"����T��?� W��ўW2��IX-�ѷx)��G��� (K=���r����A�oj�-{ؾ��t�E�N�NoPbuOQ�^�ם��i�y]�ꌑ�,�2#�h�������y)� {�'�=�G y!@ ry'4���PW���8�?$�9<���훅�/����ӚO�_~�S�����)Ի{�]!�w߾-+N�:^��K�@t����z��\��*M(�-�J��Z`�Olc��#��������#�kUV2}N?�� �������{�����gջ�vk\�E����MoM龟���5��qp�}Fq��jb�u7^�c��^�ƶS�y�rέ�Xٷ!X���;�#f`xb�!?��%��}g��$;��|�uP�7k���{��Gԧ��4C��߮�����n��Q��v��3�����pz{S���{�so���C.�%9�t��7�ɵ�ź��KY�;G�m���8'��5���{ӑ�ؿ|�˥��V#(
��p;ɍH�#��q�[��w�3�_�_g��ӝ��.��z[K�X��Ӵ��3��G��'�>��X�s��Iӫ2��wѰ�79M����� ,�LQ3��0��<�����A��Ҵ*ՈeF�u_)��0��� �  �����o^׳�^�յ��ײ�!}C[�u-OU��3��3WԫL���I%gs�r
� ��;
��H�8���D� y��G+'��Z5��9������ ,�:�#Q�v�� �CY��
�.Ib�e� >}RKT�H�z@#�Ͽ@� /��bN"�o��r<�?\��W6���18�Ȳ��v��|dWp�S� G��=X��1��~8oӑ��#+��b
]x?�� O^��?�:#�}��O��!�a:ǩ�Ǵ�V����[���(:�Zt���t.��FɯE��5Y_�5�,l�Br5jQ)�{K�?����[Op��hM�P�b��4�X5VZ�%k�*����U�v�)�^e
G%y��^�����[�i�A�	�:��5ͳ~'��%ȬA��ԑ�h��
�<&Z�N�,ť���t?x�3��8�����+E�Y4��~Q�3�� �JI�yz�:��>�t�Y��zi���b#�)��[���%)�
�<e��'�v'��];��z�i�� anYw�W�b�d
ZANBDW�xf'	�I^?y��BLh��,�!<t2�娩5\��[���|P�O8���C�|��)#W���@P=Z�w-������+�u�_���һ5~��#���s�`2��:3��D�M�qg�Ldd�� ��ʄo�O�0��E�PUXN4y�����Ֆttp��*�#ec���>:���������4��⦃�v�<�w��S�fk���$?�t��1�� -�V��Go��Ic
�-���K���y;���a���EP��|zc�=<��ݬ�=,���C�PO�*�"���1� �7�",�SDʒT ����hU��>�K�a���m�_VfR����������hIXI�Q�iǕ(1	+}��5��e���K���j?�������J���wbԌ�������d%	J�r��&� �c$A���|!.�|�H$߁���`��_�}�1�m_%o03G�X]�O��ܧ���1
�l���a�2�p��5	�*�����1��Q]���՘qR������ݖ�uA��Ld�I��4�-59/�K���~��jY�>N�5��j���H6��l8n�p�@h�J����a�!߁3uo�WS��ۛ���m���ԕQ�'�n��Qj�d��Oϕx;[��d��K�"wz3�xQgTt"�V�Dq�d��M ��zc h��rw�O��Z��:	��$\K�a��H�F�P�}1�vNX�*�r�\��b�����U >���H.	c3s�.�i���%3ni@�I)Jd
n 'uK7&cӴ#H/�~
PҮ��ر1V�Q]�u	&dR�;}�Hc%H�����e�(��2���G?�XOi��ؒ��5H�Ժ�"�tvf���[i�6*��(���A#�����eh��1�<�eⲋ㸤�bf�� 1u���z��m���;V&�>h�I5o�+�������v��GsE��E�[����q4It�C+O�:�*�eأ������Vݙ�� ��o�I?f�-��I$� ���퉑�PR,�*pL���_(����-�˸%�6đ�}1�&.�|9�̀dyK]1gG�i
b 4m���m���c�,�2#��f�yP��d�%�
[�]Yh~�vt�(`�b�[�Eo?+N�4�Li�!S�=Ҕ��*��pB˶�0�Ǖs�5,_�E3缦߉�8�U�zEK�q�u�`�E��57i�bPQ��Xl�˰Pr,dY�w��1�:�>L�d8��\��0�,9q^E��HL�FW�2&�{�)�'6�2%�T�	���
�T���A84��g��v�-D�V��N^C� ��y7��5�Ć;,$���1�p3�uF�Q����,I
���ȯ1�B62J᡺5/z4�9�%@� ��ز7'
X�;�D��!�ds�I��@�2�E�����̬=1�g]�ȸ�,�oh�YdI�:���4$�7G���䞘�r{=%�
3&0;]MC�*rx�9�� 1Ԙ�F��M]�-;%g���j�|��i:�(y|���`������9f.�평5u{�s3ŧ:���Q$9�p�hȰU��=�_&:������$LI�J�!rJ�<��Y�
�I���KO$�i�z]M��7)�Y��r�v,`�V�0ʈ:����\;µ��� C*��|�e ����z�V�E���I�T)$�j��i�$���������tԳ��)�R+b�pٖ5���xd��&%�ϓ��<,;1���>��C,�\-3œ\�ҳ�!��ǵ�21�f��ޥX�ww�gF3�������P��4����i�[d���L�0ă�+�%S e9O쟕&����s�G�t����,E�Y�:88��ʚ�5?`,r�+"�hT+�ל2s���.L�8�x�&w�L�6F�țL��.�V��~'u�Gx�$��rD����ee<�+)���`A� ��*��:�IVH��e#�T�$Fw؏��?j��:c�?����MFX�/�.[7Y���<�f�p���2�4_�G�­D��7���V����<�R<C�G{����q��D��	9���	C���;'T��t��K�oE�W�K��?���A��*J�Ɔ��ԐD�L��}=�{���uOnz�G�q5|�{M<>@���X���G�G�����Y���(�)�>��׶v����pkZ�{Nc-g��(G|R/��L�"�A�ѯ�)����SF���[Kw����+������\�!?D��	���g��~���t|�}�\��� T��[�`Ye���=!/h�+kZepډc�L�f4�^<��O�v?Q�-oancK�qS���ǰ:2wF����p��J�Q�x�V�������;�o��yv��.ז�S%9�x�h�o����F~Jz9ُw��=�~����ޱ�=�a}�v�y5�{�+���t��s����GX�fv��N�����3t܉�M6`�['���o���t�w����E �/�1O.��i��$�ĳ�I&ӮVi�hd)!A<�I��2E�߇ϋN�uk������s��%�mON�"1I-O/lw`e��ȱ�h&VQ��� �m� T�������'d�}�:n�����΍鎩��<<<u������7L���$W
٭��A6 ���j��֍Z+O��4�`�Q�}�F��Y�Q�H�IfyQ]�<�9<�K�XԵ�CQ^����(# %�j��;g�Y�%뎖�����w\���� ����~��tΕ-k��n���1��zW�Zs�=�:d��=1�E��N��g�x��-�i��,I�n��a��;-6����h�4��Gi̭%�;b
]Q��f��T~ �ݹmCy7�����T�<��k-Ǫ�c��fi�N�hѣR����k��W�������^�F���}��z�R�};�����ճr�ul���zvA����R�v���]zK"m=KS�
>�:�˾�i�>ׯc�}-����J�5�F��PG���G�b@�ݕ:���a�W�Ly��nk�w�ͨW�[����b�<si4��#M1�<]��[�Uj��:��,�Q%Q�m�N����Ou��;�����ڹlm7�:�L������ܡ��e��2bOT�q�g�:�OH莜O�FlL�jYжg� ���m��w-~�`~�t_f潩�������#X��q������G޻�_}o���bd=ԇ��}�f!:Bx�|b��L�g��bo��rԺNݖ�� �s�W�$�psu����N�׽��Ѳg|-�?q���n����E�p�_I4�i>P�uʶ�MҞ���ڟ��{(>;�����phԋ:�^����ޟ�f������A[]����>��S�WUr�m1V	>�o�6]��CCN�`����7�}��O���tM�x���4��Oun{�ҽG���^��y랙Դ�792N:����F��q��lq��<5��'ĵN����]>�l�J���چ�0YmOfG�^ċ$7d�3���|_D�F��_�}
�z{����>���U(*X�Aa�a^�t�*ح���/<3�,O+�!2����ѻ���Mgz֭����I�Q�p{å����t�4}V��G����F���u1Vڥ�8$��/L��ǆ�|.t]�d�N���W�c�z%�բ��z݉o�����hS���2��v�X�&-��?:?�t���h��[rY�,�­x��˴�� �{2�P,%ӾV�@ߎ��+��>���� z��w8���&��ҽ����>��tI��]��>������^����x�9'5��������������c�[�H�Z0O�j-�ں={ob� C�k����7��Ņ�A�7X`�4�>�����̑Jֆś�����Y���>���Y����H��
�o]��?��p��fgv:� ����Ի1��k�kN����)0p�N� {z���Au����>RN�.Y�\�l�`dFQ�έ|9k�\�#�m;rV�W��}��[�9t��ͩ-H�N�,��~��k	k��k4�ćn:A�z��mx4��M]�Z�b�]f�Ԩ��7�V�HѵTW���f���x㑆N�Cۏ`�����a���'vz��������➡m?I�pul�M�[�.��4��]ۼa�i)|�&�.���<22FM坹�^��1Y�{�T��4if�Z�>��H�'Z�����ՎB[�L%~�7�z��ω��6؃Q�Q��f���n=8�ff��#~�F%���M�����_Jv�/�=�꟨��s�����f��Ik�f��ٖ�F��T~gn{��Ug�1�c���Kw*�?�_�9ߚ�MOOۍ��� ��Ή�W��	xEh/�(T֚f�ƾ6�Gp8~��X�O�ۑ&Ⱬ�-M�MWњ֛$LK#��+U�$7+�;���!	۞���om���>���=��7p����ө��~�뮙�=����-�eOP��R��B� JC��N�͏����h� ����	uC���ӨW�v��[B��O</�kח�c[���uJ��;i�%h�y�h�Pg�b8�)t���H���Σ�b�E�-�=��Ŋ(��^]*Շ�.C3$@���L6����n�k��`u���r�}���u��_/J��x=��b�}�~��13+�`�h�^��;D�ӭ�+G�gVx�'+'��e:[�Ų��h:ǻ�|{�����ӊ��˃��0�B$�;j��嘪2�z�w����־� ж��_Z�#�JԚ��^6}@�P]��%`�<��O�b�(˲��z#�ױ~����?�V`��V�N��V�N܍W�/V�.3OV��^`�`�i��r�|Wz��&�D�ƲU0��;G�W�ڷ��1�!Z�����ҙi%=V5H��e�'Ư�xe~2R������z��G׵��؎6�F�"����li���Oj�|���6B���]�����N�dK�.��%{��m���΅�z��������Wv���oQ]O;S_�֣Id�Z���T�,S�5�:qS��G��{U����$��sX�K�i�����U��SW��P��Ox�Wy�e� E�q�KZ�ol�B������ϧКAWM���-V�$�44��������Z��X��{.�?����s������kږ����L���Vf���OU���?��o�����0ѿ&�8�����\�E���/.��Ǣt����������n�i��~6E��f�Yd��A)��9G��6\^��Ǽ����6ϻ������W�=yY՞~�p�+<H��0y��2�/8k�u��C�w�>��W������c��u6��~��It�n59i����.��zf�ަ�|:�D�~�4����"�k�U�VM���]ǡ�l���sJ�Q��)ܱ!��h��ц��Ir߼iGC� �$���4(�����۪�uTD�r�c��Q8�Q�Pސ)���y�Cعtm�請Q��a�jU�}Yݞ����~��[�ik>��n��Ǡ��+P�ٺ�X������Y��4N���\O���JډT[�c��b:��^�Y-,�"F��ɧ�Zh\Rn%b0�����tIn�����Vdc�Y"W]S�	]$�>~ܶ�G��5�����~�k����� e��C['�;�틣��kF�BW���Ut�_be��]O躅��xe'�ޘz�e��t��C�{~����ϫ�)�@���:�!�j���b`�G��喜j�Ǹ��o~�|P�Y��kiz�|� X�Y��3��ʳY�vW�V>&�0�%�=�2;��ju_�_cݎ�l�'��'���~����=w�XS3�q�z�;3.��z��0�ӤmN��b)�KhX%ۏ��L���w�V��Ԛ]��q|����#����!�R�"�|���w0�c#�3dt���;�*�kF3�TbmB��9U2'�s.��z����O�.��.��'gz�A������5���4��c(E��=]�zc�j�S�������)5��i.��H�	-	%��;O>�rE��_����� �ʞ*7��I�x/�tA�?K ;�`@�/r��F�<wl�}�{��p����Su߹��j�n�ڮ����Z?Xi�?�t�ұ���;���ҽ(��4�=j�Q�Ŏ.6�I�F�h��ֵi�ޥ�ͦF��X�i������ܒk�*Y������$���=ItZ����I�Dv�Vs��;@b8䯸� r�w��c
z�Ƌ�]>f�۝���-�3$��<�C'#Y��5����e�6��o^A��i_��'�O���|���d�F��X�"�����= 8` �8�3P�������`�؞'��� �ǯ��>� �=�~y� _��y�!��}*������9}F\y���7� � c�z��s,~�r=� ��� ��~�=���\z��ؤ����.��jY��%pk�����V��[��vn���I��U
������P�u��T���ÆpG�������R:�����;�=O'��>�����]�%��G���ó=�����H=g��:y����Q<lI/W��|YduQC� �3�[�Œ�.����k�e�%8i�w�^�O} U\�e��c$��<g���ai�UI*�z^y!��� ���J��]ǜ�22@����%������z�X�Y]Z5�S��� �����"#w���� \�瑡9�P�-���h��"!$�@o����� w�ױF��IW����y��%!T����� ��,�K�6T�jvS�QgW򀇓�v!A���?�?����dVSVE#��=� �����l���F�G'�������W��2a�tjjjf�&>��?{r���~���q��(.��4v�w����\��o�g�ԇk@&�$s��G�� ��̯ҝ1��>ZΜt�R�P�j^�v�\*�+�����c���G���h�3�pO�s�������G����$B!�������� >������|�\l��u�س�m3K�g��B���-��-����Y{����\D���s���8�?�׿��������ط"L@.���?x��ǿ~�_Uz3H�5L�.wO�>��l=}��mk��UZkS�ְ�3x4r[�r���m�S�HҚ=cOp�XF�NX�PI�>�<p��2�UK:�W��ߧ��ʠ�z���Gf|��y�8݋�� i�_����oN{m�U킚�Ieu�r{u�ھ���^6���]����n��2-*鏝�`Mk������P�Oz�+�m;J�v��Y��\� �x8
��Y
��H���H����P���� S���F�vşՍ����K�ϒz��2B��V@@[ �]��3�/���It���q>��R����ln��۰݆��n�{j�Ӵ�N���辚�0[P�����^����^N)���^]�t��o���k�z���?���m�;:�Լ��wZ��ے��'��~(cY�8�-]�fg��b�kFݻk@ݻ����Zff�lCJ����A׆4�S�'�$�y���UX���w;i�{�y>�:'�:���������{��_���_C�s��z2�I�#���7X�Ƶ���1��1����QLeb�t�<i�:������t��qҿ�k�,O�Fү�����ۊ���jDQ9I��[�����ǽSٱ�sE�{��G��f��J�y��k�dXZ}9ߋT/��/|�ٖT�`�V�N������i=��|z�}��|.��f�?�� �ݝ����4�GJ��.��\�m�8�K�����k:�3a���F�y/`�/t�s귴��ҽ)�i�VwW�j76���*�S=��^ku�u�1Ȏ#����աi�]�ۿuH?iA�n<T#Թ�V�*�~�7�V�4~�"H�A�W{zO�=��U�-��{]�V�N^_Ct7R_��Ծn�}3��g�=a\����Rkw����~�L�Nj!�o���n��� �;+@�oTѧ��ڎ_��u��*�j�I�2���&���h��P/j�+H���� J��Y�Α����5����-�k��<R��z����ʓZ�r��ʋ��]-�w��{���0�������j%�>����Htt��98'?�p鉧SQL��O3듏��&�p-��s�K���>���.��,��4.S�d]TG�3��6^3 �2?�k�ކ �=����7@�6�ۺ���O_Eܚv4�t��3(Z�a��/�>��eY�f2�m _ԏ� �Λ���;�ws"0=4hk&����+�����}3M�Ժ��?'�C$�o!������|�6�y���g�W�9�k�@�ތ�� v�F#oC��o��uRU��6���e�q�G�@6������ ����M'�7��v�����g��r��������[tΧ���!��-����zzWV�Ida����r��jI�%y�����l��goԥb-�K�b�G��CV'�̑�*�|��,1������7j�E�:{�]ѶV��X��bĶg���[[eMQ<��~��JD�C�����ٮ�w��}�{�?�_x�׺K�FWo:U�����k��x�����-c7N�:�0���3�b"�4�ڽF1s"��m���m���~ߩR��$�)�D�%���s�[/[��W��L��� $,����v�����X����<�`ם��1���@YRi QZU��da�8{���N����{����
x9]����Q�~���I�Н��u#~��R����"2���cz���#b��L��[OD�D�̷օ�a쵪H�-��5�Q	~��?�L�U]׿w�%m���zG���7/ͧH�앦i$5W���4���c�bλ{���v� ���o�n����+H�VH���x�kw�B�[k/���O\U��'���s�lJ��d��'<����:��^���mi!��k�E�Ub?�aVH&��Tx[�x��h� ;��7K���K�o����k����$Vd��~I��V�9`oRƞ38ew[���܏|]G�/q����Ѻon�eҝ/�[��{�lN���K���-=;F��V㟄qÑyB�9a0��j_Ǭ�	�z��nJu��;�2�XV?)%y,1p&�z�U��//$����'��{�h��[�F�$�uX��BNo/���E	C�*Y���~���ٸ�)![��w+��9��7н���Sy�:۵]1��ַV�����a���TmK��q٨^�5w4�톯�m-�~�k�6���u=J�C�����O����>���s��n��[����m}b��v�Q�`�IU���Z�"b�2�
y�Y��{>���b���~��.��%���ŵ��tMau޹.��Ӻs#P�ŞSg�K��x�򡛜��n&2B׆�|en����ѪmM⫥ç�Nc
�L��I�E�@k��a�r(D�<2�z~v�퓶5W�I�h˩M"��(u8Ex�\����3y{�>2�RY�����z~�v�F���'C��ZֿӴ�������}#����^6v�ԊS�հ1i�����]����ѩRZ�Ia�+'O%��=��21T%�ܐ�ǎ8����g�H�H����GERO5�^Gj��?�������;���?�B����N������]1�����؆B�~��<I�|�7M_Nd(�[dD:��������]9�������*��9x��@�(Z��n�V�$�n8�P<�s�#��#���*��p���!주��Oj���}{��f�h=5�-�}��sּe3u�,o's���`髛���Ӄb����	��܉/<���I$*�+��}� Fo��ϼ��x�v����sjH��B���� =g'pǸ�|]���t���z��ܽK#��\�M�lx����?N��&�zn��	��i��#� �� �P=����s�"_@�� �?�9����g�/c]���G�����_��>����ҙ������cc��c�j��ϯ���Ƣ�n\'�i���x�,��i�v��if?-i)hvb�]I���<�������� �U�g<� ���������{=��� ��.������f��}:XI�ZoSgj9w�y�CF�z릞ͪt��[ܠ����,|t�u����&�D~z'��c�g�{�3�>'>��`~����6�<LX ��?z�w�W��A����M�۳^�;K�u����zC�=�v�j�'S����s;S��r�ΐ���������ɢ�&..�-�X82[��y�O^ƚ�� ;���[��Cd�ץ�#� _YMkh�3�ծ�+2#Y� h� h������x����[�^����A�k=���l�^���_R׺�����#X�e�����Vx8�����L1��Y����B�o<�4�� )`9
��E�'�׸�̆��^�FƩ������bO�ۖ�� f�t�M��*�@5V�e����-�a@�l�É�l��x�XY;A��� ����؜�"�}��� ��G���j�9�t��j+?���v`+6�Yvā��VK�熺G��?����#�� W��G��?瞅r%w��nߏ�L`r%^;��.��^?���ɉ'׮���K�%f��� �=q��� ,��j���a����=~�� �j����6n\���N��DK�15��dWڌJ o���7i�XQ��yDK�@V�\�� �#�v�p|ۤr~�H�c��?O������*���Ga�E��oۗh:k��o�1��w�z{�5}g�ק4Ý�����k�u��R�CH�01����A}뒶��{klɼ�F��u]>�T�j_�^+<
ȉKLzK��|��d�C�v���Σ��6��ɲ���ٺ~��^[z��5e/dN��[��z����yMM5!���!��j�+�"�I��폸7��o����n�S'$��bC�{i���J��d�L8�E.t~x=C�ھ�Z���Az�-}-��ߍ���#w���|����E<m��Eh:ƣE$�H����)�Yӧ�2��F��Jq�N;�ݮ� ���p_r=��:J��W@t�Lh�A\���]&Z&m�]B�5�ɞ�r�~>;�
㚧��K������+�ޖ�P�=K�I=��J$�\�ވ�S牸<��%⣪�:֨�n�	�i���\�z�Fxy�K
��C$!`qܧ�=�%��Wt�Zi�S��C;���<X<5<f�7'�����2��j*�	~���(�[v�U�mݡϣ]��g�z��lG��'n�@�m��-��]$k;7_�[��V6�Y��#�Y����� ���μ1�I���Q��XˉJ��g
ܘ�R	�N�M�q �bY��hj�-<jqr�jb�	N�ފKn��
�,�r=1�)$��ނ"A͙J�m鏶;S�u�� pR�� �_&KM�mUe�C��S�K��l�%���r}1�W�\+�J�Y*� p&p��ɢ����!��P��}1��>�WW�_	&��%���A^d���a�U`B�a���5���|�7ʒ���׌yf'�BqQ錓G��d�UVq�g"�e24w�y3��	�	�T�B�2*H�-�F�Id�O܈DHJY�	%~�[v ����>Sy5 |Eek��wNafgu��vf�.�J��X藓ZMo��sQFh�+9��=��Ur�Sm��-�-B��f�*Y�=�����jh�E>A��WuU<���2j|3w�xٌ�+�� ?@��Z���mV�أ��@� b�*��'^S�s5�M˿:c���
���;M���?�o���!�)�� �pEK،@� NMT�/Y0F�4e.�I�aı�� 92Z5]�"�@���~�I��8q'�0��տl�,`&�����*�\|9�)⬸�$�,t�*�f<X�Laa�l��6H]�-%y[2̼m��	��$�m��I�t³��f�3�X�U%�)ř��b���w��8�#�2m�ҁf����������a�����ZѲ|���2(��6y�zV�Y7���+l��}�1����b|��Eb��2Ί<K��͉cA�Q�Cn�c|h�+�6�Uf�H�f�X�Z�L�� vR��<y3��������Z���y��S�N��.�Y�^JG0�<�q�&u�,O�-|L�0&�!_�7,�N���ܘ��hF��΀�4��#�����x|#������Q���*�9-�s0�
�-ŖO
��<��*�G]�zcVh�l�T4�y�����+�[���`�"��+�������͹� '����� �Lf:�nS��9+��v�5s�9oe%7U�|�'�0t��!��ր�v�Ŀ��M8;3��<����[o$�
Ǫ�q�Ns�^�沐�l0�Ñ���&��Klyzc�2���S�֎��1I�;Gt6�5dW���*hQB���U�2F_*=y?�&)Qy�6Wx/�	ĭ[w��c5i�ߔ�kƲUJ�=� !����W���ʯGौ"��n�-\R��O+�]Ip�[f��	U��u~,�Nz*�F=s�EO+4�Ɯ٧ty�	��X�y���J���`,�t;*x��?�����M�Y����[nAX��R
�qY^@�A"�G��3�I�~S����تyD�e�>@��ɔY�P���Ɍ��aɘ���OՌ_�^���nS^��w�5���U7C�hV�,��6���GU+j5���=�tU��/6\��m��X�/
�D��O�y�:60��ޡ�����,d�O�fକ3,dg�U��wZl��yww"g�B ��G�H�F�>8��$��U�q�#bv��8U,�(��ǎ������W�p��lC&˲���.����/����&�	�<���Jc� �d�r��U�,0�/��GwG�%��s��܆m�*�7ݹ;���a�p�����7,�J4�xrNw��Sm���^��2>CJC�;7D���~1�T�^-v�6,�����i��h���x�U�&Ѵ��Wg�������@mݛ�oLf&�^�i:�;]d���50���[�t�y)���������wc4O�^�%�h����4�)��� ������>+%��7#�&��I����=wO��#P�<��9U��ur�j���*����.�^C.Jd)��f�uoo�m7%��
��b�\�r�M`�������bHR�2�3����m��g��k���=�Iq�2��h�^�eW?���ո��$6P*�GvWW�z�6~���S:��Ԛ���B�IZ����o�̤r H�x�C�0���ݟԝ��E�R�.yK5%#����U�}�0��	��ϣ�b��mz�'C�{� �t7S6`�&f�H�Ljy=#����ɦfS-��5���/��`I�ط���aT�{ؠQZI�ӻ'�⍗e��Z�G��c�o\j����j!��m��G���"��q�n^�h�����*/��5d�.�����]�t�oUh}���s�Z��zץr��,|�E*:�E�F��*�D
66p��:�ʷS!�[�}iZ�=��w��U�U�V�qb�-��X-׵Z�PCE懽A!_��ϧ�4�z%������u=k�Y>n��ӳ�9�V�K�Rf�2����)'X���\:"��W�>���I��3��:/�2�y�r��	��<�s
Y|c�#Ùڭ�˹�Ar�V��1X�}�Z�'�3��Τ���pI���z�SWfܻ�Y�V����˩n�J�S�ɸL/ ���  �}�r=�w��:kS�t�i:[Jè�G�]/�v�I�jѩ��c�i���X�`�WS̃���o^T9�����0�7V����a��ړQ�� >���j�O'��x�y�YW��^���ۭ��h����tk}�jz-8t԰��������[s�=n�>��=������[Z힟�q��D�/n^�u��������������Ӵ��h�YZvm�>�/?+F���d>����·��X�xA_q6���O��q��.=��d�J���oܺ���V�0L��[+kE���uMSE����.�mm���0�յ��,�0�L�A<pMj�&St���O.��αӝ��E���Ͻ�|�z/Ot6��ߧ4���Wl.��C��`��t���������ab�@<����ƌ���m�;�[nI$�[#��cQ����HΦĽ�����SZ�����kS]G��_�n�}#��a�/�iz; I�U�q)�*¬a8T�ɻa��g��m�>��{j�z#��c}W���oC��\�4��.A�ދ�n��Ⱦ�%%�Ȝ���8ՖF$��5��P�u�XEr�H���C
��H�W��(Or�gi���]���5V���lE�*x���rIdEu*Z�2�� ��~�Go�[=������f�}�{�������;���Tc�#�����v�_Yy�Ǟ6Q������VKuȟ��{��w���l��R���C]f�	]��.mD�X�w���#�z/'�D�/��/M�5��ص^<�=�2<� L�՘�(�5V+^o!���/qP�A�]������+��G�tz�m�v�Z�FF�֝��o'��}2_5�f�h ����Z>O�ֺ��/����΍�4�g������U��S��f%��ZW��F(Ⱥ���֍+�H�rk���]�+X�c��#w������(D�N��F�;�������{�О���O��ى��O�:C���^��:冀=2�����E���C�ybc���&�C,�)�M~:� ��z��="5Gn,��0h��ũOk#�*id�ڞ�=l�� ��=ki[�SUZ��O��Չxf�/J/l@�i#{�\gm#�~���竿R���B��puM9z7���֘�"�WJiz~.����7H>���p�խ'������k9���k�B�Ezu��Gz׏��t�*]QႴ7l�$�$V���yYW>dP<��3Gt^��k��E�֝�v~�Ҿ��f�ڿ5*�$	,���C8�dt��^NUBʊ�z�ڞ�tO�����aԚdz;U�}#�:� ����j��;���y����z=1ޝ���z{���L�
��GR�;dI�j���Q6�t�n��u�
Y>j���:M��1G*���8�	&_���eT�9���Z;:���d����7pU��jZ�
�NH�>��HW��N�`yT~d,L����L�h�z?�r}�����Ը[�]��>�;O�fek�ף��w?FL���G�S�ʢ�jw�l`#E�&4��K�Q���Ž��+��~�(�jY�o�x�8m�;��5y ����e�s���� 6�{�J���p��Q�ZY�je@/�LԌ�b�� =��97��w��o��������+�ً�t���w�M�}'�X�\��}9�/T��1�!p���sh3 Ǫ��>�m��^�|�5����J3iWe�&�u ��󳈃y��a7�%U�1���8*���}����2ރ��ޣ}5->����1e���� ��B��g[e�dvh�p�	��U��ʹ�_s'���;��5}/\�-ѽ)�������V�u����o����O�'$&.���9ڐ����/~GsA��š��x�}�ޒ��<F��&�{�xD``gݱ�L�-��Q�߲��%���mh����j�qj�I��̭$�Ԫ��# �V�s{��_���Q��g���u�t4���<��ޮ�y��>Ӻ߫����Y��-�j���l�^g#'L���eu8�
A�:}�M��.�GOܣk�t��D�>j�����톟؁�"׸Шn;"��M��6vɫ�6mݶlD�ë�+R�j-[<KRP�"-bܩQ3Ȅ�����}���P�}=۟�o���j�3Н�Ҳu��N.�����t���Y�GQɞ-�S�^�x�x��gw�X���ƕ6��=W^�"Y�u-C���X�4qGV^N�������#3��;�{��;R��5�O�h$�i�e&^�^	��i�N�{-�2v�P#�QUtگ_{O�;ҹ	�>�u߸������K�y���Op]��ӭ����tu�E��� a�_������A�P|5�˭Z/[4��sW�4h���ۼW�!�^z��K��CH��r#.�*����f��Y�]����^��b���]5�ڊ���W�OQXŚ��*���!u&7O6k�:��]�қ��n��{w�̚N����ӟ�t��t�V`�O�wðx�^E��Xi���q^x���7�_	�-M�-N��:g�u���F�G����qmCE��g[#��į$��0i�):��Ik=1������c�F"�����{%=��RP���Q����~���{?�����Ns�Z%�:W���Wq4ޤ���P�Ov��]NX]'Q�VP��������M�<�d�ܝ�:������>�#wآL�<ao���j$~Z^�)����<h�hغuޠ�t����yU/,��	�J��Z)]W�r"�h�ƨ9n-w��}���zv��{�~����Ӣ�>���Vn���O�:�I5�z6c�2i'?6�9|34��2gF�ɤP�Y����K�u���_������P���apBD���UNg�6���:dwEӿbR�������I ���34�G,KI�x�om��z�������_������uvp�:Q���tWKt_�[��랹�l2:E���ٱ�_6�;� �Qɹ�Z�
/[�t�iR9U�9�P� hʱ%#���Ps��k@�y'3��;�^��Ԓзk{���{� e8�K�=���oJ{}���{:�P�W_w7M̟d�+]�eL*۴�9�Vx=a���!�y:} dY�&����A� �׽�� �/$�ʤ'	�VW��t�FP7S>�?�W�W�X~����[V�����vGQ��L�O]���B�ڞ���󕝙�fU�f�ߓ�,��&�����������v��d��� ~\Y�WuQ���'�_�?��3�R�b'������H�a�6#� ��� }��� �Qpy#�� O�� ,�]H9cG��S���b� ���^����~�܏��`Jdc��tȃ��������T�H�?_f��Y�Õa��� ,�MUVY)E[�<HR�<ٷ� ����]_�!� ���e:T��� �e�_0��+J�R�FUk�e�����t<�6Ϛ�i�E'29̥9y-n��<꽄�o~��?^��|���?L����$�T���?P<r?��w9�����LvÜW���o;8W�� � ��	���j����1v�~I�}�>�q�� �*��f�sEڨ?,x������ X��&N+-�ʁ7�t<όf����7�s��y/V�>]K/���8�����3ZZý� ן�� �=v����L?��-_�;�<��>ۮ�0 ���?��o�B[���v�x�|�9ߟgT�A>� W��8� \�q����+n���nq��',b)�KcG����6�$nW���Ļt�V��f�����x<qϠ?ϟ��ZlZ�-$�h8=���<�����=H➭9zn����Gz�`�B��Y����Y�`��
Or��b�PH����~�о[O���E/o\��2�x<}��zʚ�E�隡kh��2��v�}���}�go�ݻ�����+�ݘ�w�s��z�B�gs:����ܽ/�q�~�b��GM��c���213�H���j8�?�j�W_{�������j����a+�dy�X)��$����ԇ�.ŤدNMVBc�lG��'*+�<�k`���1W���������צ}�k��}����������B�au���-KP�Nw���Ot~N.��]=�}��5:.��9����5U�LZ��e�1!�]�UvW��M4��F�ⱪ�`�梛O��h$���m,e��R(�y#��i*42�H0�&������h�B=:�ʴ���"�X$��%�,��U��8B��m����?�/K{����<�?|���p[��;��� ��K�j����G,�g��q�o�jy��Jx��SL�t|�V�h�v)�����ZU��v��۲$�E�X+�g*a����2�� �{
�2����%���J�r����};���u/���#�f��~�%�1�9�Tuc�U�KQ�~��Ox����l{'�w��:ng[W�;;��S�z73GIo;K��uf��~��m;��H���&���΢��o���N���~�4�Z�����S��E[���玝��X7�4'�Y�y��<�d ��zgQ����>�ҝ'UJ��-� �L�e��mR�M��$��+���@�(��}����n�{��>�w��uܮ������N�vN��g!�l�Q��f}��ĺ��X*f�bî��w�Q���`�z:�W�z/��#�:�R4��.�Ҭ�:5���f����!,n;�Q��B�S���|���H�wwCꍎ�o]h^�Crݓ��ɩW�8i�k���ip�[.������Yd�3��Ǽ���������܎���N�j���yz���e�^����Zt�Pj�ffE3�d�
Ϗ�=U�|"�Od�}��ո�&��oQ�LEᆝ]*=:[������$H�d�e���ߓ�M�|!�f��V��[�v7yѻ#��<��h��3�X`�s���W����� ��7����U���vG��{B�f����к_�:�.�k�E�Y�e�L�ָ;�~$q����n>E��z�ӝ��ϋ~��۷��9�si�%��rW�TF�̭�4L��!�ʐL$X¯��n��;���{Ϥ��uڃD����U3G+�3<мhgY#f*�c�hj�2��N����1�w�Ӱ^�{�ԙ���mW;X��4��^�:6���N�Ә�����jٸI�� W7^����pG��>��~��ܝ��4�å@�����#�x��Oߴ��B�g(�b~�y�#1����Z�����F��5���ie��K2�y��D�L� ���$N���識�گ���i��Dv�Q����]ё��v����p4�<cah�[��_D�H05L��F���ϳ�XV�&wt���O�{[�Y�R��J�E�U�^䀿h�8�p<��B�Y;X�gc��çN��Z.�V�
���Wf���Y�;�)��n�y1�gt"����c�=3�K�_Idv��z� ���w�S���P��֧��tN�,��:W\t~��-#�}:�����15�uҨ�~���GQz�j=aؚ�{�M��"�w�S���I�J��E6)Y��Y�tyج��0� �-?�{�F��o��mk�'kK�F��X���3|���~ا^�h_�<Hݙ��/Y�Cܟ�.�`���3�����w[�t}�4�����]29�ˑ���n�)�Ӷڳ�)��Xkx���)뇕�$�5��v��ٻ��Mv<c��4�2W���KҲ'�&c(�g|����UY"��fA���ݛ�k��-�crt���˗�
���ķ_�3X�h^T*�F�1ߝd�]�;ߗ��� cvo��,\m�6~��t.'k=�dwOD�OJeh������#Nͦ�v�8�Q��4q�iD��n�N�uI����і�	�G%�nܚ�q2�G'�NOlq��x�K��]���I���c�dC̑Cj���+�J�@�T �;$I����x�G��{�ٞ�:��=ޮ������� �=O��}q�=OP��K����'�)<��ʏP�jX˧�Z6����Zs�9-ԟ�	u�٠nh��j�LiNH�hF�j|�,�b�����@��;5I9�7`��xѴ-Wnͷj�ٻ5I�zJڰZ�x8���� ������Շ*r:����k�����|��ب��I��ޓ�Zun����OQ���S\�ΤԲp��6X�`��NV����zm�f6j��ٻ[ln����l��"t��Py�x�Y�h$i � e����
gPNkL;[�ɶRMùv���4�5(�B4bn՝�#X�S<$�g%�$����K� Z=�?]d�_�Z�]5�h���}-Н9���n��L��d��R��=O,�Ѵ�,���͕M>���Ⱥ�~�����[^ii�@���+��̳۝����;��cU ����Yl�n�N�-)a�O��Ol5��EQ(��T�1㐠)�l?P��b�Gh;�����u�_rS��k�m3�zv�/�y�F���qk\���u}*떏��e@�(U��r��6�8i�'�E2{��"�nV@
r�ݮ	<:�0Iuk\�5֞D�����F�ހ+�dBG r������d>�F��0;����z����\��hXY�=X�M[T����]2�^��V8���t��V�gu� �0�o���+^���D;�`�BP�d�髿?d<�B61�kߏP���m'��{z��>�bh��y���ۜN�w���R��ۧot������J��պ|4��w�Q�:p����^���ӺU���btޅ<m�)O;Z��f���&�^~�����ܯ��s��H���/�>R��#�pH�#���q�����>�?O��{ǶWW�p�M�ۤ���� \b��:y'O4����:u�X����t��ud����If�֮�I���W���� ��=�K�F�$�@���s��ϩ� h���]�n�k=��f��ݫ����.����]��VO��#W��it�U��M;�n�~�q��U|��'���{Y��7`����,����p꾹VB8a��޺��)x��D�Kp�7ؖSʃ�<�n��<�����G��G���ح7T���l�}s�4��:�S��6��}>�^mz}+�p3��Q&u<�#|�
ңΉ�_}ء$ioN�������H9��>H$������I��mA$5��BU�N=�C�YQG�r@�=��]���Ǣ��Pu�N�}۾*u�S�=g�m#�:�\�Əu��C�L��f��;��j���ƌ�l�?_����6b�ӊU"H߱��9�XՏ��#*�����<�ʹ!���-ؕ������G�
�������g8�����w�����y}Q������GҴ�p�f��b�����6>)"�1{Y�Wgk[2�9���9����� �9|�/�!����O��?��dj9Y]58&b����y��ɉb
�7S���l��n ��ןc�_��y����~~���� \��7<��<|V�jH�q�V+��N ��~Wv��S����g�3?��s����?���㌮X��/�=����� �m�X��F�	�f5���"��f� ��ݏ����G��2�p	����/���w���ɩB�]�5�u�q��#�� ��;��k�9��]Z���|	��6�F /,���%�� �;(�ɕ`��#.Cq�������3	�k[4&@���G�����֎��濢��[�S3�s1���-?+"ʎ�E�?�eZ'1P��B>}d11�2!�n�x?f��P��_���f<�U�`CpÕ�����z�?_�Ϭ���'Jt���d�U�t����{B1�:J�o�B��\�ٔ��z��Z�t��60:[
�U�<�������{V��%?g�o�6O:]nMR�v�̳G���P��G�TuZ+�������M���[�ϧUI����nɎM@��2	jI�1��A������W��p2t�Q�8Ϣ�B�4�c��h����t=,�
ܝ2sWd���P�oUmU��26�7%��v�y���F��� ?�Ys�Ѿ�궴뻃��.٩���
�*F#��S��z�n}������X�������� �wGI�<mYݳX����:�O��ze>���|�gY��b�^��&tR�~���T��gK�ؚ/p����S�N"&p�J"�xGu�{���>�N�mɧ�$sQ՚��-�.IV�� 3*ב*G$�@�8�3�����1�5����ҳ�Fa��c=���$RA�'VB�fn=mf�ڛszi2�[�F�\�l{h�@�[�Dޤ�U�̰�H��mM��n�S[�:��V� Ik9�������7 <s+�� �C�.�/Vw��zZ����3�	T|~���m��?�/|��hFE�͏f�V$�"G5:��ٶ���rt�iڝ�b[@��ӋS�����L��)��N�X#Вf�z�ѯ�=ոhR���<�iՕT.ᡤߓM����1�o�R=���Z��0��'4��+�˟����vZI2���񷉒�����2���P�ԵB���V���ǶH�F�D?�# ß�<p�ڒ=��T�V�hnR���X�,l7��RA��G�O� ��8�Ni��\k/�Q�Uf~'��!@�n	��g>���
��d3_�kL�+���TKMf�v*Ē�y<Wf1�1�$��f���+�e�?����f������bC&��:7Z�&?;��W�hf���0�����;1�1V5o5�:��H͚��*ٓ���
��	�7�c)�=�HXUژ��j*�<�b�E���MYT��X����Pb�BВ<��ŦV����`J���T� ?E��*��Z���ř�1�-�5\J�	^ۄ��錦��m������5�ۃ�����%�U(	`\>��µ���l� 4�4j}�u�LJ0w^|�r[����y�d�Q2�"��_/��HA�-��QU�c"���U�q�#͸Ͳ&I�q ;Pl� i�9�2[�%��vp��:�I@�%1\��߈cU�.@e��5މ�SGna�X㉘���q��r�	?_�J��굃ĔV��V��@7��iJE������zc$c.XLm����z-h��+hx�f�@���p�Te݌�'��Α�ϑ����N,�C���s�R��0!�GU�P�|�y�"��fD�T8�J�O� sq���E��[�r�KT��U�X�Jv��a��v!����(Ҹ܀K�d�Dd1����76n(���/�c5|{4��<����h�EMIk�p*��8��	�1]�*�YW�Wh�c���8��*�R@g>J( +� ��B��JЭ�!`�(܃��Oۉݏ%p�d��{�U$�y�-�h�%y��w���;����`�M�CRV`ѥcRT���ɋ���!��,߀�F��8��oI�2�nR���F�96�8�"_o c'aη����o�Q���o�Lf:�3R��7)��ȓ ��Q������e� �O �6c��\��� �4X����P��Q���L�%��#^)e�Z��Dځ�Ff��~��G�H���5+iE��ǲ�(c�S��cj�\㨤��E�C`HL`X���z�%��Yg9I�Tv��Y �B�8m��a'�;^_�#�q)3�I][���n%��������W³>NE�t��_0VƮUj�YJW`̻Nl�CΔ�5�� ��4�&�'6t�RK�Z<��.I�c��;#"�Oܷ-��;MkB�@P��?�����c���"G��Y�|�FH2Gvh, ���w'��f,�Bo�˵Y�4���G�㻳7��x� !$V>��:����� �'c:�ՠ���
�~7�b��H��)�Ug��(�H~5^�u�9K��
|u?ء��m�f1�E�ZI���`���$Q~�GN"�5�bU��!��p� ��9�tTJ�QӒ.��I���(�K3��ʇ��0�D[�d`hbϐrE#�P�2��O.���g�����=��"���Q�u�Ԭ�UG�K%C �[���1�>2(�:�gI��nq��-�V�$R�� �?��pU�r���cek+�-(b�䓭��>BS��H��!ͨYH,`��e-����Rs���<q�Ue���I���̀�Y����W
�2�U5y�S!E������#L?�(�����@."H���FR�9�i�p���y���f
�f������;6k�*�m�1`�1�D����-H���GX���'�t����6^?�4����y14�$υ�eE � ��f�w'�N�����-�cg�Ʈ,�x�y��!Ź�M�0䫰c9��� hQ�����5����Iciv4˳��.��D�G��EfT��� x3��������æ���²wO�L���a;�KNW�ea$-|i� ���}���~]1�te����E��`��Awڋ�]� �C��ЎA�8�<���>��{��l1�):�7���G�s+���-�=��fҧ&s*lJyeZ!�,ہ�1�ίj#ӡ�����+ ��߬��+Zp��?�����cxFA�� �z~��m��Q�e�]�/&�vN��

UY��֪����?�>������ t�h[[[�9���][#;QU�\�t
�����նtG_ �n��=��� �l}mu�G����r�;�@` =�U/	��e=���vػ�o��V�&�~�J��i��UR�+ga��V?�c�-�}��=�5瓑y-1��9���@%��J�����e��<w��=l���*�X�Q_�dn���E� �y�j��8�Y�q*Y"C/o�h��Swq��d�R�\��޳�]��N����߳]�H�~��M�O�KXՉ�Ӵ}_�}1�t��L�h��?Tt�Pi�o!��*�����ޥ�Z���Z�n��K[�fn�Bޯ#�K�R�}l}$��z��[W��qϋ:Y�����$:��i⭵w���hi�����b��Kz�� �i�P�b�R�.F	(cȟ�����{y��/v������������GZ��kP�DuLt^~�^������ T�m3�G\��K|}J=Mw\���G4j�����<t5�JčF{rkڠ��#�i�Vh���C��T��Qۊ��W6N�[J�-æ��P�y,	�̒�-
�rI���J��M��v(~y���6����gt�r;�7���q���o=�]k=7�z�/����K��׵�눡����5ܪ�DE�S&X��]}*�;[��P=v�2���%��Gf1��"��$���p[�毩_�it	�ZΦc��
F ��B#"��C�뒣��L���>���u�X��d�]>��t��E�Mv���4���WZ�讌ԡ\�<��??WF7�}&�o��S�_�-���%���(Sy��o^�h��`��Z`�r�`T3�c*�w�g�^��zDھ�qh�Z2v���A����U����#8�f?N ��Gd{��g���{3��UuWQfjz�6���>�����}O%�K��"+L��&���ʭ��˻�� O6��٫->�EJ���J�H�P^Ie*JƪX�cG����Uޖ����|��Ny�,�j�)s$��(������"�vU=2����OK�i��?c���t�SmO��/q�C��:�V�<y��_%%6m���ָ����d��^M3U��8Sdׅ�}�i"�w�W�����9��>:���ܺD�]{�܍\��R��X�~9*#��q����� j^�3�_o��{���ν�{Q�2{���]��:ס�������ih��d�@�r1���|zR����U�;��zu�s�Ԯ�n4׶��%�U�y��_�,ȒA,դI㐴Kb)I�B����t�'ot3Fn��[I]��tJ����$������ۯ�b�Y^#�2�-yYx-���ftl�C�g~���q��w���V_�c�4�^��N�4��u7I��4�I�1U��E������ɬe�H�ö��4�7�Uu�t�e�@��-\�|p�04��~
��y$`}*�q����_J��}Kbtθ�w���d��d����α�;��%�{��Mڍ��=�u�hqW�z}��R�G�/k�O^k6�/�j;�YvӪ�������N@2�fRw�MW��Ft�z�3{l�v�����:�B�Z��B�v�m�n@K�e��Z^�ݚN��4u'ah/WX�Cs�;�:E�&��9V�W�W����4(���pg��{q�G[�F�����q�{m6����vN��j�KN�4�MG;�5l������^.6��b�Rj�bjX���x�K�u��ۮ��.�3�"�<zL֥Hc��H�%)f�E$���b'J֒	{`zi��tJ��֧�^*�Н&WI������%Rd�K�W��8��x��2H	8�����G���{C��n���]�L]/���Y�k��KI�џ��f�l'�t&��ivϞS���.�
x6Ts��á��㚾�IlEz[���W�3�M*�7Y'�8#�dpG=�[��lu�t�ږD�n�6*GNz��v�>n(�y&Y;̭a�eRZ5�	�t/�of]�������:Jau7SjS{a��ӻ���4��]¶�cfkp�受�������TQ}Wo������n}#I����HS�Դu(��h,W�:�Y�mwi��U��G�~���kP�{:ַ���qL�2�f���Or�Zһی�=�����6�w���zG������_@u�JufM;��m�U�V���H�4�������F�0���dTt�||�ꕞ}�̆_X���1��J�q�$��T�e����jZk�/{�u^)�����ID
Z�����z'�R�����Z��Z�6u���w�d�Z��&���1I�)Q��W@I^U�����u����ϲJ{O�o�Mw�}i֝��3�^����k:�F6�L��ɱ�M>s&����L�&�O�O�ծ���I�6��
ݕi����O���b{S��V�#�����su[⳩��ui�6��O�7V�9�Z[����>3n�5���"��L�b ��1��~���4�o'��>�zǵ9���jZ���h4wW�𖝻�|�+S��d��������/x�hss��d0��K�.�K�mZqУ��wQ�%�w�#�]��ojh����ViV�2�̓��[O���{�qwQ�z�VDw��V�*�OH8o��Q,e���?td
ל����;i����-X�1�z���ԚWVfc�k��]����zOF�\��Qt�e�iភ��!��s�9��qW�hI^�"���Z4��|�䇽Yx<���d�t��;Q��Y�a)R9�xYO�Ą;;�ke{���B��}��:�>��J���o�Y�:=�+����Ɔ"t�j{[Ԗ�~����i���[h��rg�����>�����j>�μ��$����"��'��>��ŧ8~,�42�7`dE(�B���������1�K�c[���>��^�׺�9����z�p�k����c�q����Yg�B��^p��B�?]���<2�X}
Kq�I����}p ��9|J_��s̬�����G��z?sϿ�'5''�����5v�LM��Q��͛<�,��+7�bYD��ע��V�*���,;����\�\�>�s�}�����y�y��+��c�<���G�� �c~��!]6����Qo�V�d�)�+/�O�)Q��H;|oMkH��n&D�~��H���ڟ����]㒴��X���?n��~���iީ���p1ɕ�r�[�� ����?���w��7��2�Ǉ<\� �1�QȜd���6�o���� �� >���=~O���O���<IP���#��>~�� �ׇ0�Aϳ�#6OPa\|j�W�b�A�D�G�8��3��l�?���a�>�� \���}���C��~G�fR�W'XҰ#��4����2�iFY��h������!�?P�qA���4�,C��'oq#�O����?�*j�� T�x��A>��~�h�h��K��#��\Hβ�UT�'���v�G6�5��^3�~��À��eR߆�1N�>�x� �?���d���v��f��ᳺN٢R~g����
���^?#55���U8������8���7#�Lq+c��G�z�� ��-#�__�4�#<z6>,���y��k[�� ,I����7��$�����*�
8�������	�*��^�$��֒`��n��>��px�pr���h��rֱ4����b�gbV;�(�Uk�I�#B-W�ΨZl�7Q��ҍ7Y�-����`<(��c�F �W���l��|�O�m(�e#��ξٔ�@(>�'� �'���.�����ʿ��x���Nh��t����NWk�����,l����u�b�:��^�(�.�V�Nv<�U�:[����T���ݝCJ���J��3'k��>�΅�� ��e$�^�4Cg@ѪV��G���+(b����#�ѸYX �qٮ�����wj������/h�7���{���o���%{��Q�����Z׹z��Ԗ����h�x������d�tv�D�����g�zg��'M6R�{�]�rzrk:�[y��Z��E�����������!�U�볺�  *@տi�sLݺ�I�A�W�G�V�o\$᥅�Y�-���`���!P�������r��h��:k�������j_�a��?�:gG�}����3_D�ԺW�T�����_����to��z�'T�-Nv��W&x�)�V���]���Zf��w����kK��{t�P�VBִ-X��B�x����)	{F��ڟC��7n�z泤��$6d�MSO�fX�?�o��nS�x��u����� Q��:�~\=��'A~������]%�����eٞ�uG�~���_#��Eخ��񛦻���(uL���ұF`�a���������	u������G�zm��oG��֓BӂVlj�bf��`Q�i��7=��:����F���;�K�e�1��e4�A��+�5ҕ��I��� $*�yK?��� �l�=��/�r}݌��{��̬ނ���n��Oux5�C2]m�ü�9xٝu�O�h	g�'�=JA��iZ>`����^�z��`�
�"�MBJ��z���x4J����P���E�"����wA+.]�c�H:�O�\=Vcjj�y�$F�ց�=C�v�����GR�	N�V:��~�=�����܏{�F��i�����K������u_B�#K��}kE鎰���]?]�����>=�.3���p�މ-�;��uu]��qժo�����L��:-�.8���^�q9Q �Y��ȅ�߭����nn��yv��Ѣ��V����m4�؆˙by"!�)Bw�R뚞��o�.�ԟ�4>��ɨwgG�r����+��ENN����-W�ӕs1�9y!�ڧ���>��>��i�Yg�1��"i9=���ϵg�c�sP���кj��{�oa�1⍣�T}O���90���W�7��oe�)��W�R}�v� Z������#B����M�O��:�#�1uN�H�.SL��2raLlXg�a�CO���� [�����{��Kg���^��|�n�Y3Op�xk��(D��� y#I �ڿ���޸7��v]�Z�z�]�Yu%�+Fa֯QȎK �R"��"'���:�ه�	�^�4Ί�}Ҟ����t�u�pz/#?� Ms�]'U��Kf�xzct�XI�h��#
��'�a���5�M�~�|S��ӫ��j���@�V�mu4��ȓ8�w0b���Z�F9���Y>�>��?L{�sEF=>�Ya��'/�f�6�fC�G���/��������=;���Q�>��N��W@�ޣ�Ŝ�;����98�i��G1t���ۆ.�B�=4����554���O+���N��T����A'/����Vi(��s��׎��R]?ko���^Qj�S�4��8������,����1`�ٱ>��+7�/�� ��{Y����K�ơ���\��պCM�����FfͲoX�ڎ���؍�ؚ#�ii�k�o����~��zu�6��+P�b�:j�5��:Obyj~�J���FĒ�iة&�|�����V�����wu��ֱgP	5�Q�]^
Ћ\��ܺG3�E�bN��F�ob�_���O@���f��N����d/uGg5n�ei����ǿI��:ޚ�^���3�Y���l�a�`�E*�E�n�oMGR�hgt����rמw�$��c�&�EI��Dxe2�h�YI��^�l�3G��&�5)U�k�J剂����w)�8�YSĬx}��ө{S�u��d�o]��:[�:�7�=O�i��^��~��3���vi�qc�+�wM+_��48(��4�c�w&�ؚv�Q��e��1j��4��eQ:����;��8e����rQ��m����=�[H�b�Zk4ɡ�Y"����yC�}nOmT�ߧGY��ۏn��{��y�ٞ�z_Q����U��T�E�5��|:�W�˦�����	���d��1�&�j>hJj��F�WO��+�z�-7C�Ri:�E�&��V��e��x���K�����O�n_�;�|i6�k��]E��<��lҊV�#ȡd�w���A�kj^�������>�v�H�>]>Ǭ�E���Cк3L���tWR�	���V3��w������}��,g���JS�[mJ��_�uk���D"gde'��#�`�B�{G�� ��k�04�"�7���X*�{~�\{�d�[�8��K�ga���WC�������z-�m1��b�Z&�����v�5ܥ/��:�V���|L�l���MriIH��k�%7��B���b@��^�!�����p	T$:n�%�z�@l*X�}��c�NO\|��9*=g����n��� x:�W�^�����K�!��n��Z"v�0#�cV���3�tcG�n���BŘ�����xh/��e�-���/,E�+4D�:8>7��{�~�Ȉ���^����AQ�z=�pV2�Xp\�=zOG��9i��� w������Z�g.�L�>�t~�M�=��Τ���ݷ�L
�:Q�,R����V�ٙ��ד̠߲�I<��X�O?v$� 豅@��= >Á�z���3��� I^��ܞ���3��]�k�8y�'��'�]E�f@���������ݼ�`�֦�$Mfѝ<ρ�aoJ:f��7�w��W�
�X/<q�G��|�v�-;w�ХI��>܎�	�<����{�����tWFk>�{��Y=��E�����O��C�Zn4���v~��2Jر��,z�������ʗ��R����� iT�[1�yS���xKZ����J���<]ߤ���\� 2}{{�3��=��_�s�ׯ�-�vϣ���u^�wp"�#��Η������MWx����_��	X%|��	���Ȫo�&�
���#�~�H�2����x����M��v����IH=�}#��@|���䏿�2�y���#��w_o��ZuN��`��ڧ}uMR�~�? �-�g�Zx���G���2H�P��ղ.�9h�?b���ڝ�$���D�9#�Y��<����>�A ���4t+Uݡ%�$�O �\@�G�G���R`����J[&´���JW.�t�����gޙ�l��������~V4�%9r����G$���{��ȣ����s����� �WPɶ�洿'��`�6~%Ib6(?��c��z�{i�d������̇��:�IzaV��LI���4�n\����>������WdV��Q����~G�~���+ {;'��9���g���%�2ru��f�����x���,�l�d��sn � ����X�������G?c��~��5��!+(����q�� �
�I�	��3K��vǭ�mL{�0�x��ݗ%qorFİ���G�R^%z���R
�P=}�����뤟=�ag`���8-�>����;��V���:뢱����?X��I�>,�r�q2�5Z��2牌t���`�����jkGMI,i���N�B!��>ԀG�G�@� #2�Bk��ۨ�'�#N@���s���>��n�O�b�O��O�����_�zK�n���u7p-���H�.?o�c�FҺ�����z�M��}���O���j�~-���U�*;ų�z�ۆ޽��vεR���O	�j�>Ck��'��H?ڡ�{h��Q�}Oݺ�H5Y�۷#���2�k9���cY����1P��OJ���A��;�=w�/k}��wm���ƛ��wL������=7V�wYuL��n��M�q4�l���U��'N�R�.�ݣd�Pu���ugQ�����n��5Y֫C�,J���e�G�@�)Q�Z���:��5���]�/�Ħ²�~Gq$����)Zw����F� d�?!l�]~]q����=W��L�OX�C]��;��i���S��]�8���ű�[�P��;}���_���oz1�wtj���7�����hf�[�� �%_�?c��������7�ܚ����	�H���%��Ĕ'����M}z�c��_�{�c��W3��z�1tmDҥ-7��}?�:kC�H��~G.g�]����%��mm���s�Ť�4k����K��x��=�����|�O�@����:��e�5KV�N�}�D�9 �Ӷ8���F���$��^�t��t����{������ײ�˸];�i]:5��2��s��[�z=F�{�W��U�U�a}_�5��ҭ�_���Z��Z���>�R���ڎ�إ��%X�!���!��ѝ���^�l۝a�6�m��Hjte����j�8��A���<2/����_uS��i�s=�hoWvT�m#����{o�t�z'NZ� ^���΁ZK(��/(���Y(�����]t�����WM�#���QOZ�#����3��s�H����f��m�BƧyjK���{	(n9O�	"#����Gp�Կ�C^��p���;3��u�mw�v�н��2z�D��ȶ��E/���j�_k6��ȫ���l���'��2Ӻ��mr�Yj����xF����Ԥx[�R���E�>9D^(myk<�R]�$�#���t���n�C�]׵��΋�7 Y��y�Z ZA�6�*�-|FY<b%�zğ^��|�����_����>��HuF�Ӻ�I�Q�i��ȱ�%�>Kc�P�D�����-Y�i�7��~"��]�e�c�n�Ih�}�O\�Ix� �6'��Y�tү���Lw�Vh���{�-E�H_� ���{�e �\��E�I-Q1#�!nn��ۍ�{�I(�A��ܡ�<�G�rc��03�C\���6�`h(13v���V�7&o�b������L1�2B���,��e �4��>�C.J�Y7��	��I��јE�NG~S��oVR�<��/����1�rX	#*M|-B��X͸��G�m�7�r����+>����Ȼ�j�$�y3�l)�+Wi�
���J�d���Zj*C0�,|(o���-�g��8`�#������Lc��l�]x��t���6G1PށX�Pq�4�
�!i�T~F��@�76B�!٘�Z|��1����Ճ�yh�/�myQ|�����Ñ!	Wm�c�/	S 1<��%[��ʁ�>_$+�+5��d�dB�f�Z�x(n8�(�.R�7�O�y��-ɸ�X����$�q�)i����B�U��أ-�Y��c��/�4�;�edEA�
��L����	a��^�A����QUj���I&�,>�Rj�N�yzc#��%3:o�2IM ����m�#��b9����%�J��Jh����F]�ZM?�|�o�EZ���QX��uK�-�i$WQ���$w�ͫ���l�wc()o=�3?*�R2p��S�A��m7fo!V�M�匤F2�&�Y�OY��Wp*UD*dy�6��N.	c�d�$�AP��x����2��})�V �#�A݌,@�O���+A��]����i�]��~ ��
r��ȓ%�*��(�R����+�@3dƆ;I���5�ԩ���N����wuT
X+�'u`^X�D�Z�#�'ˑ\e����2��'R]�d����ɋ�J�M �*8�˂;}vC��#m�6Lf&�2]<�I�,B�ʀ�ݐ*�U�D�lQ�پą���E�Uoz�	��<\�7-�G�<#f	�+�TE��^I3T��%�9��k��E 0��rT3�$�c6a� A�/�|�W�<����T�Ϧ1�V��ZU'zY1j��5ѓ�	Hso�aĲ�W��1��"U��4��Ej�#4
�Ȟ'�>X,�&���c;y���gM�e"M%���tv��?�,ד0V1�f�aR|ժƶ�.��a�J��s-��,dt6'"�J�D�Y��U���Ϛ�ʫ�qE�QSrX�MҹUz�jS�_%���(̢��݋~ߌ��"�O錐��<r����ȟ�V�u�+�"�B*�y_���������m<�ȮS��"N2a��H(��;��Q��c�,�(bV�j=��LX"8�֫����}���1�(2�U����:QA������w`	B�쳟��L�y����D&���?�T�SUW���|��"�µn� �E^4Ȇ<[�H6j��Yf��l��36��ǉ&z��J_eBNUr�������ys@�PW�+錓yR��j�q5y���gQ�ۓ?� ���7>YX�
m��ST��2IK� �1���N��Z���P�ʭHo$�+D5�$�*,�)6y~3!uG�S�Hmبe^V����(�8R�[��wI@/������o�'f0`������Ry
��tf'�,��<����YUvٌ.ʫ4V�:;33�����T|���3Z�� ;o����>Ӎ Y6W}��Č�����4@M��أ7�K?O�2��H��^�����0̨���HP}��Vb\�Y��mս�j��G����e�,�+� Y]ef��D���<y4c4��^�0s���J�����<qe�_L_�=�,ק�rd
q�p;RE��/z������|\ҙyѡ[���}E�gL�LBRb��j�|G��]��������iu�|�CF#s4� �"�d��5�)�+	$���ur��-�~��ї�ad7�Y2�X���;��*��e��pŝY@��>C�ȭ��iƩ�j5u}P�K��7tS��$C� ��������L�z�N��軛I���-*����I�b���h%_�x�ʟh�Fᑕ�9�]��Lz:ڱ�^�i��c��w;%u.�P�h��q���|��7?�y�4`We�Μ�Bh��VѺ�*��_���8�%;��-��iHO�2�Un}��y���}om=��ѠۗFfK�nK�n�C2Ą-��}�[�{�5����Α�ǸΒ�r4�ܜ�C��΋��y�&e�.�e� *���6F8�`�uh�,��k}S�]-�,�Z��v��Y^;5�eV�u��Y[� �AǶgG�Yt[{�&��4�zҡ��J�Ug[t�*�Y��!�P��Q�!�b:�	���E�K���C�?m��OK�>����b骍<}3X״�RZ�m��d�N3"9��|P��?�G�Jͫ�5��:������c��<R�~I��� ��@�+��o�g����	!޻Z��F��眈��,w��H���v�wA�D�`���V����o}�v�u�G�/X�#��Z���/N��`���T�G�yt�E��A��HP��^��T���q���!y9�s�D:��W1K��I:�淨L�� ��E���2=��k=��R� T\?�晛�ۗw��&�=CK��mf������j|���.i���@�;�9�s�8�8Z��i���P٭�����K6=G�����1�Z� ��mmwZ�'g�S�̿��H}��X�k6�X�$R9쐌̞��.�������+�7@k���|z-z;M�OV]M�t����_7���+1�?)��R�.HǬ�M�^�O��T��4ޓn��u�/bQBE�[���=o<i9���Y`r�7|m"3�g��wO���uKA�}��!��j�ۥ�����QVq�9�h�c�oȨ�Z;=��g���r]e��t�Zh�3�:7^��7l4���v��3I�o��i]u���SfOR�c���1�d�T8F�Qy��/��=����i�͍>c�ȓC��Z{RxcGf�M��	����������^��,-}sM����Fc�x�xKv���0B,3G�D!�����6�{A������=��f��=��_[�izWF�Gw5�t��m/�p�iz�&��d�de�+3S���omv�m�m�Ս��ٳ4��k�d���M3Or
L5g�#Xz�y�8���PL��D��ݝ�� ���Q4�ڻR�j�h�u%{W ��Z��8Y�����+?o9���O�#�<u�c�t�|�	���tG]ug���m�hz�f#�c�?/
�R��o!�͍L��Qǖ��n����'��]�GuO4w4�}Abj�'������y �P�,h��q��-�~w����;f�yj���r�[-6Q�Kd�,�K$�q"������~�ÿ�����u���q�c�΃hk�����u:��Z�HK�N:�� v���i�������[�7z��n8��kN�ef�I娮r���������m"S�iG�^�c��� IWK�m����+����nb&T��k����3���� ͛�n���?�'����#�Gv���Y�v��|�=P��m"zF^7�L��K#5l�q��U�!ԍ����:��/���o���:��Yԥk:�N�W�R[1'��=���ĊbD��� �>"TH�Ӯ��To'�;R{{/Cҡ���Ig�&J��$��谫J�Y�_���/�ǡ]�����%tx�Ow{-�>�v��ߪ�������jZFF����`�������Z4�c_P����<oʆ�.��Ԛ[�L���az�7u�$z<ڒߡ�*K�A�d����!��Wr���2)������t���a{��m#�j�Nu)k,o�n�é��.��*�/ă������~������;���֝����f/Pv�x�C헹����]GQ�?V�j\��]GS|����*�k�>;�|b&�_Zn�ݗj��M#P�35���JլVc/��j�9,�rHݙĄ�w7�6���}+��Ѹ6��+�t܈,k�e��ư��ڬ	���ճr��t��|���?r�m�MO��X:.�ތq������ �p�7�]#��Ki�A���L�/ ����lYLc����KV��ק�R��ͺ�s%���T��t�X�W��$O �1�ߑJ�]��]���K�kR�	I�/��s���B�;'�Uh��O�9ɾ�2}�{��t�/����Ovi��x�[��������f4L�,}K�{���cW[�M�f�~�G'�'�����M����&���j[dR�q�(`�`Ӗ�T,C9(ihӟq��E��" �@�=�z�A5���f��j��">�cS����ٍCG�Z�H�֐v�)�~����_���^�|���_���� �izˠ;�ӽw��)�u��������gu�6q�龮�a����t��K��5W
3U�u��������ƃgq҂ܪ{d�rQ+"_�a>�>X<I$���",�B��z���ݧ^7[�X�kj2��fd���D$����I�����F�HKI
��牾տP�u��4��V��� A�^���O�����n��zCQ�4�S=��4��?�Q��i��Ӳi$ka�sq��؎�)�vHa�"���a#P�cD��D�l3yT��P_�. k2U�%Ev��E ���KHиd�7'�T,��b��o������^��:������.��Mc���|�L<<k3&�Ӛ^&J�hF&F�xr��X�V���C�2��Tz+���A� ��Ϡ��q������x$q����G��I$眖�Q��|J� ���#֖6����[bd���Rvn� ��m���3[z�Oi��I P;���oל��m���-\U~J0�ԓ�~�������Z��F=Q������Ȭ�v�4Z;�Fp�� ������*��)t#�
;Gi�O������ؿ���M%��\7w?P#��8�~ǟ��.}w���<L�%�|���}.T���3�&��`o��m�m��YV�4�ZY�vS�x>B;W���'�y ���,z�Ũ=t���h���yc�� C�� 3\����Xd_E8v.��u?�$ϋ�����`C���䶗u�}��?�P�T���9�3%��vZ�П�����䏿���i�eūb�A�p�w(�7o�m� ��[G!P�e>�ehd�.G�9�Γ�ӌ�A5��I5%�%Ӟۡ�j�0��Y>(�����8Hy}� /�� �9�����=s���=�?�f��KT��W���óO~+%ʌl�T��b4M��R=\�U����~��� /���#eQXr;��� ��sd�����WH�L�N��� �������j#%*P�4h(c�4_��q���f2ƕ��<�����nG����
�HBvz }�y�� _�����i왚ff���J._;Yx|2SrQ_u|�To�Ğ �������Ub�ZK�I�0KpI��8�}���M"m]��*ֆ?}�@�`~�������Y�iZ�����ZGSW_"q��7��e[V��S����������G���r��!<�����=���}�����m߇�zs��"� %���~�� v�ۧq{����=�쮵��n�VWU���8i����jz���un�Բ'�}.�5lD���|�C'K��N�j���K���"��*���#��NX�J����P�����tk;T���6�l�W�R��F�1ɝc�D�'o��;��طQC�����.�u�Dw�z�W�>��~����������A���v��z��/Ed[P����/��2sk.��5]4]d��F��6����[�d�pj"�Y�wjR��=*��Z�Դ�'�P�yZq����#��Z��ꦽ��}6�:a�$���P�V���Υ)�%�HyU�U��#ֵZHI�:��=A����;�{� �p4N���s�:?�n��%z��q�[Z�|\]���g\�V[���Tê�VjwQ���d�i�Ĕq�F�73[�\>('[�U7$���8�Q'�uh֥0�@��#^Px2��$9���_�in�t.VI��K�ty���K���� Y%-#?tva��HU�3%u�o�#�,l�f1��ۯr=��ߌ��@{2�s��;��5���%��e�X�t��v�4W�ci��i}G���-O+)1qYn����eub?��w>��m���l�M"�u�ԓ�ů�q���5��Y���ў�y�F'��g�]9�s��}
��M	G�J�3���~jϥj����n�*j0Cj������������>�{o�.��Z�o\�>ǻQ�eu�j�8:aS�r���Ws�i%�Y�j�����x�;R������a��a�i}!Ѻ�uίm��֥��i:���-+��ځ5:6�΅�]Z���U2|�k!�5�R�^��mZ���r���n�ͦW��R*��"���[/ +J�݂V	������3�r�C�~�;�]���gQ�2w������twPiz���ھ����ރ�Ա-'�#'���l�o˦��77��H��
Z���a3F�E�1���.jF����r;l�q���4��$m���OvW���2�ԝ�O��k��I�A\T��x"��s#�$�{;��O�G���U��q�_��>�v��=�t55�F����4���e���g���-���[34�d��i�+�wǆ��w��;�L�(jRQ�x��hbxeY$���`�?�Gi#�Ē�F�4�Y߽S�D܉�m�.�����D�7��I%�'��	!,<�B�)y���I8�}���{=�����oGtb��{~�?X�3��϶��
z�H�t�uNgPfj�2��//I�㧑1��8y� #a=f>�I�u��m������>Z�~ǘGe�+�'ƽ�#"�$�G�>���9���Π�Dnmfkۅ4�sH#�Z���Ig���4�zo5����C����_���Ox:��:����u�g��F�^��^�ܽgE�l����=_;U�<A�a�H�þ-���Z+,��n����5�ѫi��u�S�x'J���V&�C�+Ov�\_4���C)z��
�,�[EԗD��mJ���nM v�&���IR���$.8�?һs�G��ר�����u��~�{����H�_DG�;���iz.EOw{7G�f��m3Sӧ����!�%#H�ZV�S�v� ��"�����m�ýoG]VYӶ��u��x�iW-���Y�����,����?��wgjO�b֬ۆh+��K����-7e����t��}�Yl��	־��{�����]�p��]��q:{�uo��Nt� Ovӭ���qt�O3��<����ff���F6Ll�-S$��6�Ez/�ݽ�w~��sr�
�.GJ��Z�3�M�չ_���"��5�>�A��Z:��}Ƿ6������Wv[�����>+�H�m�t��@�F�dx����{�����'�x>�z���]hzF/I�o����r����^6��c�d�1�gt�R_*��|�S#�~-�.*��'z����7��7Qֵ��C9��.�Y#YUhU� ����B��ᔜ�OJ�zx����ҥTY�Z}{�D�#��'��=�W������e�}]e�^ܻi��oj4��{h�� p:v���&��z�6��Ώ�2:Y����/Rb>��M �F�F��$V�}?/F�[��˫j�g��m]�^G�E5Z�j�bY%�8�/$Eg�4����Q�C��X� h� ���t�H7V�;i��Z��l�3
�Z�E<�T��J��-W�#�@��!�� {������6��k�����~�z��:wA꾥�~���QҴ]cS�����@�zd5~��S�><��ҳ[aj9ɸq�zgҍ���t��ݺt3�j�Q4�FβR�aڬ��,�+��X���-{�U�m������7�QJ���+Ad`�,խ�X�@�k�� D2LG��{��C�����n��g]%��W?������������Z��=I�uF�돋���j���\윏��0r��_�D�뷨k��Y�����H{�1x�D��W� �PF�da�0�����m���6�=/@�O	�lq*F�װ��Y��ܙF�Q�$��z������g�^����G��>��22t�[����:ϩzK�'��֤F7Q�V�8�ƚWY�L:�4�-WwnCnȰ�d����Q'r}$���l���=�)+��<kkl�����vS@Fc<� *�{J��$Fh���`��������v砺jX���'Nw]Ǉm�e�Lk���ų�'�rt�v;qa���=�c�_q��!�{�����Ϋ��Y��4g�����gs����z�F�20?�Z2�ߍ�a�?ٔ `}}}C���[�����O�����ר𴌍�=��^��jڭ2d����HfU3:'�eF�L^����M�*
��H	���]�K�Z��</��Sʳzg����'��X�Ո�`�kyI��,G؏�Ea�E$~��#F;=�q>����ڮ���w�����>�����1��RڧZ�#���2i``���u�Uu*�# ���,�ۏl�¯�9>ϯ�$� !��W*BO
����G��C������5{�G�u���G�����iz��.�jzu_F�k���c�׳���q�I�j�k�%3%�
6<�1�������D�wO���7ar�>����1>�` < 	��Vw0G;Fǁʏ��ABð�������)�績���uV?p�������{Z��.����5���.^nF��j�� ^~�U�e֘z^B�>MC�(��WSyh��T�	��t)���dT�|��ǎE^9�Wغ���Z�Z����v�����I����.{�79?A��o��=���?�}1�]�oY���;��ڞ���w�q3:Ӽ�ҙ�1t��z��Y�v�>�ʞ.�������Ƀ��\�:T���^(�:r��Eu19t ����2�!��G��g���j>X坞���bp�G#�.W���ݒ'x����f������os���u�V��S����������_�����չ�����:��f�sQ���FM;o��:���E^���'o�X���?��f��Z�Y�![�>���O��c�'횑��d�J��|�F����hyҟ,��|TQ��!��&�������a������p����쟿���A�������A��6�`h�H�}A�v�C#N���<��� �Y����Oߏ|� ���X�s�54�^"\�VEe�����7#��?$� �Wl'q������>�?��2�e|`�|���ߧ��j��:$t���juP��i�4o�`N�v#}��.т|����_���_��ψmJ���w����u~n���z7:y8�d�`��Cx�H�QǓx�d$�@m��1���4֥�!��I;9�9��w�ST�:9���)���_��q34��iN��hϋ����Щ�u$퍤��
u%�LƾL��by�m���|d���(_Y_O��{�q�ى� m��p�%Y߅A��o s��l[½-'H��*1�ok7�� v�w.�y�U��@��綯f=��l��{���ܽ�{������=�w�Y���p:Aҳ��_3�{�N��O�����u�&�бuM�t�@$o�y�qk��M���cS�{m��t)�j� ohN��mF��Yb��ZH5Z�ۧ4\� |���}��j0vh��h�escbb�o2�$�K)���|3i�~^U$���������R��%�+��;��+^�^��'m:��4:[���۬a�9�K�]�D����R�>��c<,�s?V�NFRK/5������͓�t]�GsX�ږ)�u��Ѱ�<�ϪC�2С 4��^tJ�s��)�+b��KW�7y����IU��IV�&+],ڮD���Y#%f1 6چ��~�^�=���=�t/�>���F�}�'���f�5�i05��iq��}['V���i�L�W���W\\i�f*;R���֖�ӯ�:�����4-by�����8���U	c,g�*���Sv�C���I�j���{1Y�X?hi�F��f)��B�~��I���u �	��Q���+;�S��^���Eә���3Z�:� �^�ʤ8`u�?p�+��b:/�0����
�b%��V����P��[Q�4Gk^��_�;�'�m*��}U�o�X��X�j�;��D���/O��N��������u�h�L��^�����ts.�_]�?lJIU�w@����=9��ʻ��� n]�}�����~X��g*�^g\��$����Q���<��5�������r<�9c<� ��T4K�H�cY��R�ԫ�זs+.�)�H[����X���¯����L��*�Z���Mn��	��� ��%:lrK�e���d�TP<�O!�h}�w�?����WG��>�t���;ӝE�����;s����q�
h�:��\�l=��[P���L,�?��_�]�Rz�6�b�+:n�	SZ�z�i�%�0X�IT�Аq�~�|�	���]v'F�l�Lݩ�i����f�֨��֙��j4Ĳ4���G�^���鮺�5rzϦ��u}�n��u�rj�6�ܜ�;t�j���/�F��hN��|i�&s�7���Gb�ZE����uu�p@�˧���H҅��U$�U=��rx��j���S{[��[{�P��X� t��.%oJ��b�E��Yy� �v��k��Ѻ��HhX�7����,��Abwz��G�4�i�t\]CY��.�Q�jR�5[��):�l����3~��4-aº����ΐ�ZEjp�*���>����ZiG�Y�I���Co�ۓl�����=B	쵔�cMx�BWx噡��K<1�w$�;�u=�u��U�ս��QN�t_L{x�t��mO���Z��������q�Xj������la����n�j}b�7.�V�y9C�Me��W�� t�޴��$��F�.=��D�O��tb�صH�k�����i>P�	��lZD��"����;y�*�Z�q��������N�w���oq��=
�'��֯���U��җ_L
O��yc�q�q�xF���>�t����:��ݺoJ��cO�.�d��vى|�f����d��@��dg�b}q��w��[�wP؛#T��F�ԭǧ�zD�����"2V2t��8�Ʃ,
35giC�dKM�n�ꮁ��)�[@�M/���4�Y�QYk%i8�!���J��M�cqm]Km�"�5}SNc��	��	���b?J�=��X��� 9�=��*�
��(��o��J�v�z�Bŕ����I4?�&[�jk����KM�Ҋ,�rlY�đ�@X0A�̇#�b���� ������,���#�R3W�y�V,
�6��c$�U�LxW$��jw�<�goˠɼ�*�ΥN��"F��hATd�,���*�,Zf�L�6�ߛW`�o�D�c���˒�U���#����0�Au�S�ͱ�z�#�NL����[cqǛK�O�֒�@�eIR���r�/���g_iC�3t�����_U �-m�1Q�vO*P�
��nTQ�)\�oDm������o�M�e<�t)*
ZyNQ7����6�����wWQ���I�õvS�(�ez	$���F����ŷ��f1�����Z���Ql�����x�����v^ ��v0�S��C��!�p��G�Dݝ�z��)��qܱ���|����D����E��<iP���`��؆�c�9����B��*&證&(��h�,7 �%Rޘ�,����ezq�8��h�"21�b��0��^w�Ɣ-;=_ű�Lڄ� �9)Ww"'��zc(ͪX�ZXЕLr��P�_#+����ܢ*��1���c(�Ti�(^*$V^M�D �GA I�&��`��+I��G{QM�WRӪ�e�0�*����b}1�o���W$4�D�� ��3�3rD~$q ,@ӿ����Y�q�F9P��G|�R
��:�jC��M9}��َ���̬\�%)���� K��|d��n@)4Ȕ�����nq�4Wd�'��W����e�}��w���55}PailUC=���P .ƭɾ>O#�� '���bՖ4cx� ��͌XRB�i ��X�wnL��JX���Lc��Ҥ���z3f�ip�5-��P��9|$���\�B�ⴢ�LV ;�
/�Ǜɐ� "����V1/�Dёy�-��9���� 6,� 0⪫�Pl���M���&��z:�ĭ>w��	;#�N@>�6ǖ�`'�S%I
g9��:Όի� �[l' �x�TޘĜ<����Gr7u�'*"��A񪲹(�U�rB��4�$�0���-�0�B��l�D�ʔ�H�_�w��#�oWdRI/��]���&�Vi���y>��� �J3N-��"����W.��*�� ��y2��1�ZG"�v�����u~)uY�Xcc��f'ɀQ�w>�ø~L�Q4,/����3x�|TU`&�XQ����B}1��b$��n� �AnT|O��?Vvo��m��1w�����fD3R�y@�Y��69v���(K9e ��(�4B��!�5�rBdM�@F��M��yЀ7!��Q��b\Ib���J���F���=m�}�fgY����`���c���+�1��վ4�B�� �k�J�c@�/����
���Y�i?|��s@��<e��-�pn
ԛ<����b4���)�5�7�nm6�N�	g���c%�b���0�f�F>6�7%d��=� R�rn �pvae}�'!�zPΩ�� �H�)E�˻8gQ�0���+_�\? �L�|��2���߃l�JM�e(Co錦�Zugvo0�&ro:�K$�.�r>�̰�l�O�2��x�9Ϋu.�,���Ҧ4Y��:��۱��(��U���F�W̙I�`�1	�����"�ȳ+�؏Le3�� d�;�*��%���~@����޼�����YuK�������X@�;\H����38c���m�Ÿ��c5Ǭ;K�j��Ɔ>/�6���]<�'.��]r!U��b���l�Dn*�l�hq=�躝��ɛ�ƙ�xk5��Bp�ɒ��1��B��q ��Lg8���<��E�t����򵥙�E�V�O�h2�Լ4�D�V�C:�45,f��:Η\�J�SlJx�D�;MT����O ?�
N���W��}��u>����}C�1r��=�edWC�'�t�4-�ݗ��?�;�$�ą�����z�G�_��_M�O�{���J9��ߞ�v���2di��Y�7}�7w���H_X�-���#�j�{a��d����_��Wo���� T����M�.��f�)��N�S#������M7��������H���=]��چ���e����GӦ�!�Q�*�P(�����#���nꆱ����6��]WC�Z5�kWy����b3���X�V��P�D6f�=vf4�i�}\C��].6��3�d˞\ ��I^��_&�$�0�Y�}n>�ճ�F�w��@*���A�$���z'� ���s@�.�˹'�?O�[Ked�ېH /j�W�<)n�o\n�{��:�ޟo�5����om=����G�n=�����'A��+�a���a�O�0�pd���X���0�\�5��}~�w�ޱ���vܖwVǞGa>�-����ҽ���H��<rD/��D�G"�H�����wE6�ΏE�0W��
�+��>Ru*��i�-�5c�7hmS2ױ���Gÿ�C��δ��÷���=����᮵��<�a�ێ��֣��O�V�d�ˋ��bR3��m5<�S�0�Q]��V�f�靝��[�&��6}k�{��|�6D��Q#�6D�I#D�H@�֯���lN��Z�M�WJ����jW���b�QZhlXԬ�	5+q�*��}=��2���7�����q�j�I��蜽Nx�*�%����^�����OZ�l6D��V'����/z<ڊ�iu�v�mE�_׮Hg	�����1�Cդ�����|/w��	IuW�s� ݂s�7{������?h}�wｚ�����i���ު讴�mE�;W�Ѵ�;��2W�(&�p�����}6ڎW|��]���I���n��{��:��=�~��B��v�騺���3C:ج�a�xı�I�nI^��3|Yl��ﰺ��õ�~�J��r���VF��8�a���ee���7dUw��oZ�?�~ܻ���/\u����{������������Ӻn��ft��Ņ/��]�/Dv��NVVDgQ�|;�3~���R�_n�M�|�L<�S��R���GJ=�$��"DY�~�|P펰����C�������u��������n�֍"���F�X�T�eU���G�}ެ�����7�^��W��n�W��s��_�PbTb�7ݓ�&=Uy+�e*N����ӦէҴ��R�N�54�W� �f2���������M�����!�u�Z��;�.MT=/��'�A+\�s1��Vv7��п���Y��k��[��U��ڮ�v��ִ�cL�]j:~�Lhc�GU�}3V�1���@�@�9�����߅ؾ,l�T�Y�C|݉J��$�m�0Af)�Z��(�Q��h��A++loD�"��!�M:��*�׻5���|̶!x��^K�z)A��*����N��Z��������q�����Ovt��_�מ��c(����G�4�ccGX�rj�(���^VS�"���j�#�&��^���4)��n�4rO9��c�#�;"VeT�,��#P9_z��u{P��zyA�}׫G5:	�
u��|Ibil7|�5ʪG�Ā{�Ƿ�����jݓ�7�E�}\��LXu׵^��%�=�϶��<�Һ��&��W��̊iytR��*��� �-ߺ���lV��i��+�U(ku�ݘ�&��+K$�KX��E�6��[]���+�V��mR�N[:=��RwAfN�*Hei�q�	㑛�ս����ݬ��eս������ t�3;��݂�^I]kR����s�=��W��]J��*Z����b�s�>^V�1'Q6���J�U����!�X���D�Nx�X���b��X�XE�hgNb�Y��S*�v�Cu:56���v�׷�Y�(ݕ�ڕ��h�i	�CFB\�+J�	M%�Y�`�һ����{Y�/p���s��=�k]�}g�:�3R�3�i�vף��ϴz6�%[9b��"�c�V��m�"O��=���w%�,i�n+����y$�Od"�M\D-?s	�ͺ>-��ߚ_O�n�l�sJx��#���")���%���T#��ů���g����3�Yݓ���?�����=��d��Ϋ���N��������N���yg꙲�_��r�F��{�������mWMj�Чf/2Ʊ�E�4�� !�D�@�J�nC)��������4M��ZG��X��Z�y�Yռ��b	��,P+�3�znXs��&N2:�E�[b )\ܥ��A�o1l��)J$�j�,�v[d���x��^�g����D}�>��x��c�9��9��<�� ?��� �7Q��l\�<-9������2�lL���ݪ�+2�b[n&�������1�U���唸`x���8�Ϭ΅�#�J6�Z4�Q��<}����#j:�_�+l�C,ڦF\^�A%���$�U�$7�r]���&�Z�y\Fx�1�>�[��{�{�^�bIY��tS�����a�#�� s��ݺ�0����cgs��c�d��~I-A�=�������n z��4�~$��Z>�wq��,8oC�=��
�[����K\�c�Ĩ�����������tޝ�Þ#E�r��3.T�vg��ţ�&`�C��ďX&���3ة8�A�i_`����`�^����̋J��C�8X�R�����G���Ì��^��{������cT����sj�L�Ģ���I����RŢ@�,=|R�5�&�IV�;;[����}p@�� �>nkZj�+��Ӟyr88?�sw�����󮙬h띎~�^J����=F��?4�,�A�=_��aZ@�?����Ϧ���x�O�9�	��q���N=�_�3O�o������N�w��u����{?l}�����x�[&U���:{�u�yں���T�R�!�Nf���#N���l���u��$��3W����r��C�K,����L�x9k�_����+K���DP�%e�B�vO2����b9�OfQ�~��_pm�w��}��e�/�n���R���C��tn��u[_7Ū�/=+z���$�_k�[N/V;�5��c��&�	V<Fa��$�f�yzM�/zu���P�x'� pԺ}��t�hXRy�./�_YԱ01��cd����e�6ǘ  �f�Ay���Ɵ�ʳ^�W�.Ih��/򾛟g�Ԑr� �iv���d��1f���D�?�rs7Gis�蚆�2s�퍦K\�������P��5+3m�,�Q�ޱ���n����̒����҂O�h;�����,��^�k�mv���L�Ȅ�y@��f�Gی�o��l/�{��o��计�Gv2{c�k�%����u�I�j9��p���I�㏕�Z|�kjCD������Z�hW ��	�wF�o]������,s���J��`���
P���IZ6@A��}bۛb]=#�h���CvńjR+!d8�%�BH�#rj��ӎ���zo@h}!�D�GK�&ֺZ�:�D��:�Y[�_P�!o��M����h]��-<kT1�l}CNўXW�Si\Ƀ\����Iu]OgT�V���d+[R���Z�$�0vR�u
�)ԩ11��%j�1y�O�D���ꞟ�.����<�d���bV39�Q����Ԡ� 6�� E!����^����C�7�}k����^-��/�׶Β���_�H�L�{��K�e�i���4�/Y��KR�rs#}WE|1Y�&5���3�j=�)^�R�f�(m�KP��Kb�2�&ں��VO�H�>Z�"A�`
{���v�G|�N䯧��X�JJz�lK�i���5������g�2�����g�N�{����m�O|N��zJ�x4�w�S��H��'��&pɍ���u�{�Yyҏ<-	4�gA�!�*&\�m3�+M�>CU�6�n�2�O�h.���:�9�W��Y�a;G?[��$�� {�_�-T�:]���_�R��x��+��M��;^��'��㹎�w;�����ez�ޖ�߭{�=�c,tr������ T�I�M#L���q:7۟K�P��{B�n����}w7z�����Xd�G�=Q��sF�^��WԠ؟��\�,�M;snf��ͭ�_�\fxiVw�'�G�b�Sa^���M˷,̖u�_6�[��V&�X�sXY���,Of^�!�ns;�^�;K�t�S{��'����p{��H=���������+�umJ��.�]Q�����k����g��9j��^"g���w�:�S��d��m������%�*[0��$t~b��e��?��j	y��J���r�� ���������F��E��Eu�V��'kQC<)�+�]Z���7�T������ι�3�=]�T�L�^�GTB;�N���{u�ES.����;韍���S_ȼ�mZ����dP����e-j֡G{jմ�O�h��
y��u���G�$����� }G�L�oj�[�b�^�VeP�{���k Q´7Obp�����g{}�˲�_�������u-y;o��v/O3���S�tN��?��0_\:��<�ve��B�D���g]4O�
5�Y�j1h�U0If���ݻ���Ӫ��i>V$��<Qƞ(�D���tg��>)o>����ٚ��zk3ԣN�;ei�|�G�G7�����<�&��8��+�1�m��|�S߮��4�Kh�}��5>���uH.��s�GQ�NPkĖN)wӃ��ޑ�2ham��w��E�]]WL�e����Ѵ��&)$<V�a�}B`4,T俼��vϊ��?K�J��Z����;������L��=��r�/l��8��� RN���&G\i��������A�����9�/p]�mԕ5.���j�^#���1{�Sd5���K����4�~���k��K�k[Լf��U�J�z�p߳�;H��y�G�5Z�n��zV����nU�Ze���j���;,ҽ*������=����$��ݑ��[�Gg}����^oS{�����ҽ��ߗ�:&e�4�!6�r��	���s�ru�Ub&,�J��k��ғoR�^׵ �b��g�iWQ<��k/3�$*���=�?�n�?��7Q寭�0ܗO�����B8�-��Ս�O,��l�Һ�� #)���w����@�߹�ٻ}��}��������ֺ��:ã��#@������%gmo��Z�r���T�΢l����5�%}RmJ�5���'t`��"����	!�\��+� 	ܝ��v��i�h:\�e�����%�"���xʨ*J�q"�����?P�t]��wd{5�n����W�E��C�����ޠ�2:ST��<���v�8ϫs�"1�ަ8z��a���
������ʖ��;ϧ�Z��h/zXh�Sj4���`Y`9%�i���y�q�9Ū��~�stlM���;z�Ԗ-]VQaa��Q_R��x
��3��������.��e��=���m���{۬4���#�z��wL���b���?�fxp�&5t<i��bA�[3R-Bqb�m��:+F=��[3�v���\j�%�}�ITK�fy�r��c+���t
�hݻ�]�˶�oh��U�r*S6Zs<��du̱��x��K��3��k�t� U����t����f���}H�z[�z���L`t֛�Q�]�I�h�W�h8��S��Ѱs�o���/���>ldٞ�⌻�XӮ׸nN�Ĳ��O<N�XЖĥ;�BUO�y�@�;5�2��iU���"�aVd�X�5S�h�~�@���Y����h�H�=��;��������?V��S�?N��Q�m�I�E�!�5L���c��j��?�]�]�Lִғ�g��R�}uR$���i ��<�l��U��,]G� ��/������<��s��q���.��a�jZϼ��t�v�F:�j;{ڭ[#����M2sV���Mp&k::�fD���T�6>R^0��rʵ>t�ɮ�|SD!�	f+"����d�^�q��U�\����&v����H-�L} �� ��Y�
7a�9����Vw�,�ޙ����������G��+c+O�:�-l��]�lv�mO1�gǆ���c񀡚vvvw2H�Y���'���v��?sSJ��>�8���C���Ͼs<{�.����_r:� X�b=�����ۻ�i(�7Yj9v�Lv�H�21ӫ5j��}A�t� Mr/��8��w/��R��ʜ�����s��'� �SO^�,���އ'�O�?�����} w�ۧt��vcL�O�>�i:G�,\K�����k����"�}]�mN��Ժ�Gow�����Û���a/z�#I�ݨ�t�د̸�E��'�y��ߙ������Ԫ�Rʹ㕅HR� ���!���l�� j}��w��=/َ�ߩ�w���԰zOP�������]U�#]K�����M�ׯ�(1	���Y�;�C��g�m"(���+�?��+*8 �X� }�����S�c�J��R� ����
�D$0�`I�r~���w��.�:�Z�c��{i�+�ڎ5�ޣ�r�#��}иɐ�-3��$m+��u��Zv2`a�c�jY��W��7�%�@æ,!J��ݙ� ����~�	?� {34Ѩ�P�;��ڪB�}K����:��� <z��8y�}��7t��R���u6�սW��P�5w\��Jf8��|'	*i�Tq�9b`��س�K3A��\��2�я"���*�H
��Q��zs�� ���Pz�g��}���$���uK��IN\��`�Cri��F��ylTl��/�x���1�ݤq�ʂD��Q��<��"zK�B�����%���v�hH#��Q@���KK�3��~����?A런'�~�!t�Ow��?�eϢq���+A)��G�,��S�D�/�Tr��	;��?)V�;G�'?����8��g-�y�n�~9� ��� \�9LMN��0+z��;H/%Y�G(���ĀG��7������v�����ۏ~������<ݓ"	�~����2/�u4�3�����)1a��C8�R����)�[bO�o��#�����T��tB��<{<x����2�}=�<���3s���������][��������{���wI�֥���S�tO��~��ȋ��O�t̘�j:Xu�\�a3^�e��i������v��GC�V�[��Or�p���c��� �ȧ��7V�}�j�̓xH,��	 #��]�_�!�}����,Fw�I�o;u������zoT�������D{��k�{�쯼���9S�����M#Mӳ�[�������.���|�/��MG?&�8�_Q�D͢m�;�����ں$T5���mhR�%=}�����3���t'��k6*y*X��G�(R5��j[��}7S����jPA��5:�<�9�S���bRG��a��,�Ν���|��=��*�Ə�ǥ� N��_WtF���]C�wn}M���:[�k��=�~��
eee�N�Ƨ��?@9ƅ߂i%_����'}nN��E�$�`�,U���c!v�*��1�.yd��=���J}�4��kų�\��I��Y/�2 񏚵+��}Y;S��ʯ���}���{>���;�ԙ~�I���\�ޭ~��w�M�Щ���Qs���ct��_�s?�CN��r1��[�X�����R�{����sK��l�I�($�>�ki9H�ҡT�mg�
�_�Y�d{17!�>���Gg�ݻ�m
6oh�؞	�ArH�h�Y�� i��9��D�Ɵ{橗�����(w]~�]/خ�􇷚{��}��+Q��{�]��OA��b�k+�c�e��WItܟO��a閻�V˶f��eI�f�az�6�@5M�j�m���jP�z:4/jk�����D�b��S�EQu�*7ohLa]��}fk�Vέ�'�څ��CU���TӪ�Ȓ��,3On{�ࢰ.���c��������J�+��Oq�/��њ����k=���6���,uVj��5\�����EM�2<�U�|X[�/���m�x�J�wluU$�Z[QA`&hi�{ ��K��5iC�f����,�M�.���j���rc*�W�XUJ�&)&t�	s;����������_������zs;�?�ν�����~�>�۝_V����P�k���\KO+Qǋo���P�P�}:w�Y�w'S+j�K|i�k�NM5n������N%X�Z�4����e���P�a�n�=����[UMv�վF;�k�Y5
��H�=b�3����2���P�� �)w�︾����|;�ޮ��ͳ4�j�f��=E}33Il�'Ͻ0ie��2g���y�+��A��z���ܳb��ںF����#�(k�RN �5'����������7�Uu�joǭ�[e��I����E�w��)���`��_t�w}��0�+�M�]E�����5_�]�����j���Ŗ�*����;�'S����˵Nr��)�� �O�}���~�W�KW�Z�ƣzj�_�+4�J�B;��sAU�/�Q�\��:��#�l��j���ƇM���JJm��I��d����ZQ(u�E���ֿ�+/V��ö}��w۾���O�.���غL14�����g6�cN��\��ͳ2r�#%4���x[,��v�7Q5������Q���KRj���*��;�Xx_�T�iB����вI���_?N���v���%�oM�R=�h͆�W�X%�Z�X���bH��q F~��w�Ϊ�u����?Qt4�2%��}��:91e?,�;jS�0���$�Q̹;�]=����M�j�ߣ���d�]:+E����I�
�������:��B֧�nMG@�Jڔ��^@LA8=��
>たO+�}��?���f~��N�h�#Й}=�.�t���=?�L��O`�5L���0���������T�33�o��:���'�w��׽�����=���rId*�� �^jY�,��J�W����G$a��o�����oa�u�E2�a�wvҒ5Z�h��,K7,�OI��U~�C���w��M���Du����Mj��V.��h��t4́M$���=O��e}er'�~}p�E�*'�jP��� �~���ͻt*۷D[�t�ʚ�O-Z}#��� ��Pj,��>u�R@#��0o����-���-���ɥj,��4���|��m/���xX�#,l6ṵ�ތ�{�=5������j�=l�L�-#��E\��o����|��� �[k��VT-ɶ���+�$�U��z�3w藵�0�����Y�&�Xn3(?I��a�]�^,��|=X��{O���J��Ɍ��ni%���ZjQ��� �~y�WM��[^}#Tֲ4�L܏�Z~�u�|D�t=;_��ZU�U�''FAo٦�٫-+sR�>Zj�c��'���rb.�(̤{�y�u��j�6k�|V:`ùy�2?�T�`9�����5n���f���l�n�C�������GN��>��m+B˦�c�u6�=Z�o����luVXU2>��
:[T6T���'����2� ����N+nmf[ч�$��\�㰞�}�,��Xr~ߠ�?�߿~� wW�t^��ew��zw0�u�n��:_FȤ�.��}s�綝�i8�J�'d�
)`b��i$�E�Ą��HN� pD#���`�/��|�o$@�B��`䯌z��<���v��3����Mڮ��S�ݱ�NfS�vR:,���4;�ftv��K���W��;>�u6��=)25i��s/��Ӥ��|���Wx;D�	=�=���G���@s�}rO���@Y��Q��� �9���l��1ֵ�)HO̊������̘�!�k��C�`��(O^鏣:�Z�X(n2�����#2��c�QM�YWa�}��TK+���^6HV��ն,���1JI�T�R��9쾘�c���-5�dTBhr,R[1|i�Ѕ�.�NX��n�aQv����ߑU�e�(���n�;с]�ڌ(;zc�Z�U1�\X�<kR��1dF��� K3�y"�`@oLbv<�wR��Ș�����gT)����n�!�������!�7��2Lx[��Y�qɸ����4�9�]�4T��ʲXQC&�Y��]���F��}��c���Ɩ�8�t�M��6�O�JNZ�><W~L���`j�8Ң�P�Y1�K��3�ʯ�O:Rk�3Mw��<�1���$4	�����ey�;��Sȋ>*�a���S�)x��"T��qky1�CZ �����F,YU�Ewf(@c:�vq�̚�y����1��.;*�.�� %��9�]�����y�k�1��Y||�>���v*zc��ҳ���4σw���Y�㙧��b̿+�l1��P�H��+EW�<�¥m:���*+m��'�� ���RoE(9Ό�qJ���iEk��j ��	��Hc��>��`�ԉ�~�=�>> ����*�Y���<K!4�o-4@6����1P��S�3���PcRL�K�P��9��x��5}�(���Q��f1�)�!�AQvo*���]Ĭ��ٸ.��
1����6Y��"�\��ˁ(�P��'��d�ːR����z����)U�-�iHZS> 9#Ѕf��9�/�Lc��Q(�%DS��ec��7H���hy�ݏ$!�8�,a2�����i63���C�*�f�'��I���URG؀�G�aW��HL������4Z����G�/&�uPf2d�u�;��qQ�TPCA�gBY�O� '�c
C"���f��}E��뷛� �o3��ܵ8�8m����Fȃ� ��D����|�X��<l�@E��LbZ�Df�V/���six\�9e&���(�D��wj�0�yd⽧(�+ ��9M��+���1A�P�l ��q��W�֥��޸��H��M^�O<9�l��8 �^L�,���R��Y�1�*RrJ+1p��Zy*��~l~N�`�ˈ��9��%<��2P��\�gT�!ɛ�Z��.�g���ޘ�D�u4��.�	W�%c�*QU�/"C�#��H��v0�2�FئA�;c�"�r&P�UNC��h����>�P(v2��V(�c�8��|�p�X��_�:����a�ScSw��t�;NJ��c�K`��)���1�|kTJ�%i����L����qYF<f�N_@�P��+LeZZ8�ʹ�5G\�ij��&��W���vb�SbI=1��e�'��]��V�'���w�ʍ@�%�Ď$��0ƴ9�b�@d�$�36-����P���[f�ƭ�����[4�l�Z-�y.4����m���̀�Ōd^)��P��LM,"Zk;\���ю̠�X��yƜ�K���\m
�Ȳ�*��G$nJ� ,dk��8�Qe��Ufr?"R���}�Ѷ�0��� ���3�j�5���X��C�[!�a���T?��
��Y�i��'݋�=��^��b��){d�>>>-i[ձ�	^�."���@�Z�TS�63�^�=���*����韟�j����2����Ѩ�\@H�+�� ���Wu�e/Ӻ�ˑ|�Yd���B�����BJ�f~*�d���Tͦ�/_��~N$3
�ei��]�L��tYJ[@2��(�T��f�&׵k6)؂�KV�f��G$n>Ύ�20�2�s��j�+�R�t�R��TY"�62I�GF���?����߽n�톳��-��SE���g�����ii�q��:��IH�rF��s�?�p�5}-��P�z��22ũKۯ)F�U=Y����UOx2��uk\�k�v��~t��oj��W�E�����*Źj��B��L��h�V�^��/_�ܧl�}G�:_���Ǜb#��L��+�L�����j���T
-���J7n�������jĸ�b�ȁ�I��E�<{%NtVe���S��`�Qנ���'�O�WV�fe���l����Za��째l'��������H2W����2��xa�u���v�%��]sO�ǩ�������R�:�O��C,O���7Y~������u_�{�I�i�Gx���,j~fKb���i�L��Ff����ӳu.�uU�z�ۃb�uES�E�ԝ-�4Kr(Sʵl�<3Y�H"qH2Xd^��%��ݻ�ot����ӽ�:�Ojڶ���_����`��3p����_35��u��$�"�/�$�=�~�E�(S}V]f��>@�Y�<��*��Fk�X��v�#<����+}
�I���Zl�JĚ\^�B����Ut�('I���_h��&��$x:���'�T?q=���n�'Iv7;�v��u�q��z'G�\~��M'+��2��jzF�^P��q�mU���e�V���[I��Z������f�6����e��r���R�;ܻ��'������⻨V7����Gؕ���S�5"ЍG�;��A]�ʎ��&�أ���U�~ڽ�{��(�����{��,n��֥�j]�}a�O��M`�]p.�����F6R�b� ��9r����jL��]��%�/l��K�7a�;uk�1��������V�&��vxX$�6En.��[� �x��n�mߴ��5K�im$�+Ge�_1�4QL;dD�h�KDΌ�r���?Om���>�����U��v���NտH�u�Luuz�O��u=rh�0�j�a�['+M���l�7������('�i_KU/sX1���ظ�^��(�,
�8,⺒x�>����+{JĿ1CO�)��DWT��h�� ��?9 ��"6v�G.��]�'�=��^����;�OL�+�n��M'�=�ԧ�bj��V�������w����SΒ�� I�<��^�m�ﵾ����wy�.�n�GD�M^(�9�NR(�D��cܱ��X�v�-k�� phZ��'D��3Q�fxd��'�4�$�N�U_�^�EP��/ܫ�{m�ww��gVto�oo=�������&Vf�՚gA�M\��:n^Tc�[*9'�&Fa>���[�=2������[tG���N���n�J�o��۪�<��������Ħ&����h�7�F7��vv���U���$�.ԓO�<"7K1C�dvxEU%d�c2������?F?s=��=��7U�K��Q՚�뎻���6�Թxr��0���1rm���4$�	��,������*��?��յ*:��'����".��3����6�V���o�0�d�N���i����b��Zn�r���A��lI<K�D�¬̃���TyP�<�ν��k�S���������Ǵ�#�t��|�]m����e�s���Ӱt9�+�1�ԊefT��Z����8��J��H���PA-��x4�u"��yAwY��g��Ux���kڦ�cCy�M��]���`j���8��<0�@��'��"RO�A��n�tc��t֍����� {�a�*i�]�ޮ�OH������F&^��ҽb2�u��<�c+bk����l��#QRɶ�T��ܺ���l�Զ�k��m2�[�mC:�����8
�$�o���ﱒtZښ6���F�7%]*h�M��E�N�-��5h �) n�̡��A�_���.���`��t>��y=a���� Ҏ�w������k'G��O�;���ސ�?����G��o������c[�!�e�=Z
64]Ct��܅�zV�D� ���a�<ecw�"y�PJ�Dg̷A��ij�z�Z����X��:��>��)Z�c����{�H9�X{Q����z݇�Om�]��� X�֯�d��h�I�-OL���MqTeǆf&Z��# �a���1o,�OTz�6�P��S���5p���� ��C�0�=�&ɸ$��d��h�W���nT� s�$pA�oכP��Th���Ӟ6n2N9��eW�q�-��\s�5A� �z��潈T�*������~���	�x�G�ʋ"X�4+ܮ{������#��?��?( ұƭ���9E���.I�V���ģo��}��O�Ѱ�Ο��J2�@�
���W�Ü��v�$=���,9<����}���KN����ۻ�I�1턹�Ӥ���WVz̕n7>�a��D̱�$�� Ff�A�O�|}�-6��L;O<�pG�=fG���:q�Ժ��NѪ���k|MKR�Tz�6>.ȷU��%8�~Hy|	7nWԡ�ߴU����R�D�?����s��Y���v��ܠ7.��pps� �{����}�w�L��<v��[���O�Zv��dks�;`�晗�W'R�]L��|_�5ы�����͐�6o���FMZ��UgE���s�vPR��	zP�O�Oy��f35��x�ݪ'�S���#��{C�����R�P9ڿn�^�?MOp�/��˱=O����t}[Y�Q�=r{=�<��c�vk���[���5#�5>�'��&=?��i��#&C��wT46����U�R2��\�4����i�r�	��S�w���oT�Z�zM��:}qs�]8�a�8n$��G 	ؤ��]��@H�ӓ���ߨ_b��u� ez��)�����uh���-OQ�N���{I�}@�ջ-��u����������])�#�X�k�۷`��-�j���K�-��ç�6��V1jH�0]?��i���ۖ����J�M5kV�I^�H��e@�b�*�Oፗ�d��g��'���<�zX�֍�{�ڧ���� W�I�/r^�;}Ճ�5�GO�zs�7J��Ki_�׬[M�[[Z����V[��ec���Yb-n�����k`o�n֕����%��6�9�Y��bZ��m�� �Z��VHc >T�Y���˸66��mH�I�=Y�zP*v�m���
�C*��)h���I�d����w�}?E�u;e�]k�{y���NuD�#�ƭ���X�W�'�>�X�鮤�Qc^4��<��{Fߦ��o+�kB�g���m��
�N�$�f�mԄh�Q�4]�"s)�[�gM�c�75��hU����-�\�Ė#�#jv[��gƈ���ѐپ]��-�n��� n�w�X����t(��{��Һn;�N���m5>������7Lun^F����Miz�5n�]~�.����6�jf4��M��t�m��5�#S�:����>F���=f��v{Wf�Ԥ��]�ζe�D�ݽ�]��omm������ڌ�[�V�)�2�Պ(���%���&��p�GE~��~غ���L� k=�ӽ����FM=���g�1��v3R�5-[#X�sz��u�c�Y�{m��v�t��.�3��(��k|M�����ѓ{�ѧ�S�����U�{#	[X��x��+/i� i��	��y$
�d~��6�)k�;{W�5&���$�P��f%�S���Z}�8���w3v�PL�]�� @������g�7ܯz!��Z�K�c�E�� w}��SHӦ�g{{*5�Ϭts��荏�=;[D�%�c�,��ΐwR����!�V���Nͣ�	$�^��=���Ins-���My�6����=AkZ����콊$~���-����Y���sR�1��S�PAY{+J#KŨD�H�;���9ӱ�(n2�c���'K���>��ێ�v׶]�յ>�������t����n�qz�Z�k����_o��|�#�޿��6d��N�q3s%���t��W:�\�M��Kv�}>�����^F�t�6��*��?����Zt���g��,�G�Y7�Tkuj�wR�&�#�|F�}��۫\	��H��WilI(�ƽ�����O��Qh�����4�o�}7�tn��ogݩ�F�=�v��#�4�u]�?z��?����Z�n.P̮Sc����3y����uN�ȃuk���sRյ�5����b������W�*A4�Dy$����wn�E�ޣ�h:zy*W�i�%,� .gY죡�2��E�$�N��.���� N?�C�֓��t�_�޺�� \�tg\����_S��Z��Q�iil�n�c���r��a���;$���:O��FN��}�w`�25=Z���x��+(qW��dp�״��(�V|�v�]�������C_p�qy�\@c���a��e&�o����7o�H��`x�<e=��gp�ܯ��������3ݮ���oy;��-W�]��tG��u����:N�����K���e���x�ʻX��/�v��v�o�[�tϽ� ��/�]"���d�Dv%��c1Đ���L΁���o���֭GM�5�~]��M&�J��S�/1F���		�����{v��HOd�ɏe{������i����]3�X��Sӹ�֋-K'�:�	�3T���[M��|�?"���,��Ƈ����/k�4h&Ѵ�+J�$Z妁�>��X�M�i"D	()�2]��6�����i�����K�T�oe;ନDh�0+7zs�:�{��?�?O��t�hz+� H;��#�>���=ڎ��'H�wTj9ZF������d�l5����2�kQ��{����#�3�B��zF���E�}co�W�oM�lN�]�5,=^c��@�P�)��X�<X���!ֵ-��i�vF��?M�,�ASS���ƫb(�G�Ν���si�9o�p|�-������{M��컴��:��Th}����ŎV���A��P����5�SM���˨V��3�%V��§;�間���wݺN��C,r�%kIbͣ����d�z�H�s
�]Y���l�:yۺ��b�X�O!��.��,TE��`ǿ�㔲�Ѱ�[3w{k�P���U�۞�t��>��ǣ����N�뮖��Ώ=;��oK�j:
�u^���8xٙj�|�D�r��蚵�/�m�ku��K�>�]
�%*:mkEĳ'{i!��	#y���P���6˧{m�Sp>�SPy��w�Kv͹��fh֫�u��Xʏ"X�Sm�s�˶��{7�_|~�{��tg=�B��tި���Eu.�������K�=���ľM���x��ހ�����!u�z��d�V�[�V��[�L���W�-�2�5l
���b�y�9�����\�J2S�� f��Ƿ��{�j�m@ކ��q��S�ĒW��F�����j��j2����s���'���h������;ӽ���{��ע���qn����^5m����.W*`�a��:v�����zk�s���۷6���[�[�֕b�$����؅��$�i*J��r2�_�r�)ĶoҖ���-�V�Ơy|��X�֝?�����<k�ͯ�f��]��=�Ұ;��]	�I���սi����K��[������ӞzF� �P��X�cO4�u]U-U�����[�pO_D֬m�OgH*i�|�4㈔�aY�X�/ E#�4Q���m�t�oh�g�4*ۇT�Ue�oQ�n�nIT<ӷ�:D�;���n���7����кc����jt�D{��Gu�Nk���V��z������z{�_7�h��'�a�]�J+�VVh4o���֥zY�kS��L�]�I)fU�{9%\8�답Y�w�>�H��i�]z��i�W֫E��F��� 9	!{x� g%}���^��	�.��/h�����z������_�q:'����7F����r�Y�F���3uL\8`5)����ެ�Mb���J�X)�ȱ�#v$}A(f���~��>��˜�V��@�&+�3��G*��D�~���X���oC�?��鮏�z���t�6�z��q���{��^]G�2m��c����l�����r�����z��Y���Z���7n_�����y� ,A�� 

�t5Y�7w��� ���R�d � �{�<�[�c�Wt)�fguu���cO��j]I՝M�f�OHд�t����Ò�2IcB1M��{#�%�QG�� � = ?���9s�9���� ��{'�}gѯ�� ��3��+��ow]	�wK��n��/��ո�GL�����7��W�2?/Q�HӦq �K*�9�lyӅ,a{	4U$�����<@�����yc���~��HeC*z$�J��@���?�#�~�q������ߧ��#Z��ޖ���h����%��n�Ė��t���CF:gL�yT��^�8ʣ�Rӵ�^��,0
	R� ��:$�?c޼��@q�a:���^f2�!b� p���Q�d?��O$pߞ6��?������p�zӣ:�ۖ��=��U�Pd�=�(�?�>�A]CI�\��8��(g����l��$xn�oF�e���%y#g
='�B{d���a�P;��Q�׿�d��I)ux�	� ;]�K
y�����_�Ǧ���{���W�7Gv_����=����G�ow�3�+������:@̇�6X7���%x��tE\t��Z��8B�=����+�l}�rB�}���륿mjo#�}/�����s'o�C�S�s�X� �6l��d1#8L��AD����?��ۏ��劑E$-[�I<���瞱[�A"�o��C��L'������Tf��n�����O,�#r��}� �������(�K�$�����u�6`lz^�E�Ǒ9����o&�a�m�~���r�=�T���I���r�!����� ��y��Ϧ�;�:6�v�8d�TrFV_�c6}�����{z]x�r����~�z��g�7�X0^�H���_o�� �OMG��#�CV�PiYG�bN��|���?�Y�j:�wht���#绽;��O���֧BX��byY�ݍ�菹���m-V�-$�SѴJZ�Ե�[)/I�$�\Я-�R���� :�����uxܺ�!<qp8�}@�p>� ����,5,_�٫�Pr����s����������{����^{P�>����;s�SU�m���)�
-�O>�]�v�S� ���w4�.��ԵO����
��{�z���C[߻q��������2��Ǩ��2i��*��2�����f��6��kL�ʎ�"q��>�Z2���8�Hx��C$r)�@�ۣ�x�여;��g�mF��˫5��R�+�2�C�_w�����1���[�ZÆ���.�����4�#J��|�x�6*���>w&��]%����O���9K�e:�e��-��`�ՙ�y%�Ĳ��c�{��£��R�Vp]���G�%�H�5m��4�rxG��|G^(��I
��/�	��y}�{��?~���-�?T��a�ZƼk�u.�߯l=��#V�4]/O��c��M�rs�5\F��Ǝ��m#Y�Ȅ����HuOF�G��e:���c��^�SN�+�����ZCf��E�f�X�Z�Tf!j=����n��LF�-�2Xd$��F�+_��Hh&^�^��q��߻��.�vS]�K{�Խ�vk�]^�#�;���?H{��>�M?;M�����֍n���Ny�>n�����[/0�r��w���ΐA�����;���t��芒���x<��X)Qt�#+ g�\Sc��XT��'Rw�hڋ��wv��L���D74��9"4ƺ�S��n�>�]����'���4{=]ҽ׽}�Oo�	���f�����w���z�R��;����:Wo��@��^��4�G���,l��&�W�[g[�t�[;Q��q[��fyt��jif���Zhe#�d�XԥG�����6��%��?X�V���+V�sS�^��5��<��n�� ƒ A][@d຅�� g��}�~�~�2��wC���Niz�>�4���Jgt�P��A��>�Ո�9���e*�������Kc�`0�@�M�(���4�6��#��H�&�V�R��	��',��鼲������|7l�����]6���#N�.�ի;�!8�b9}�F�9��s��'5W�~�=�{�?v�����OU�=��Zj})јZ�n��8Q�%.xS�հr���(�ǛO�/>/�U�~���_Ӯ�l����^̯[q�j�ٸ�yk�JO�bx�ĝ���Vc�{�����S:�ѭ��v���Zڻ~�CR�>%t�ߺ'c�2(x�� �ͺ�&z�H��=w�Ϩkߞ��'@bk�����f�u��@��D�,�O�1#,X�VI��ά������#�n��t�H���Z���Q49�i���Z9�dQf^c3<�r>B� |-��F�u���� �ç׃�X��]G&�P���=���RοP�]��y���������5N��-KJ�7M�~�.���G�����Z�Zu7TE������!�#�L�<�U�wȊ/v'^7֧����v΅�Aq!q^��#����n;*��^�\�{+�:MӺ�V��۾-V��+��Zs�a�k⮵��l7*�PI�]YC�/z�Q�>�=��c���{��~��8�L�r:'�:�X����K�`&~��zf���E���'�gKD�H�� w���4��t�mn^��ά�%��a�ح�8l<�(#ʫ���w��x�;��L����nGJ�akO6��ذa�r�BK5�IUT,��A1��3�h�� Ln�ts=�t�o���:ǨkӚ�{g�w�?P�p� ���� ���uM�s���Ӧ�X���� �z_�=
���-V�P�M�� mB=!#G:x�,>Tn��A/��B~��Y��ζ���~��NZ�&�����-E�?�~�w�̵�����Jɝ^��~�zo�m�t/m��i/�di9����'hB��`�:���:�ᇍҋ4��q�MmBt��?+o>���z�6yJ�?�B�$j�!��e5$/��$yI����;���ěd[�����iË�Ȱ�b��{���I҅�����Y�{�:O�!ӽ�CWӺ�[�lG�zg��Β�g�M"�} ���[i	���TT�Q*�JT������^��X�l�ɡS�$zlڷ���#�����Ỉ��UJ�*���Wh��b��Ej]�~�/�A��ZAg�*�4t�d��uJ3���f��C��z݄��x=���:A��'z�sz[�2#�������s5z���+N�m��r<����D���u����:/�jt�u���֪%�R�N$�x�و4.'��(Oo��E�/�gEv���=o�z�T���w�e�^�vWY�T�eD��"ԙ�yaEi���L�V^�v���q��k�=�ץ��R����u.��?LtfL�0񵞠�G7�z�9K�$00�g������m�E�
q�jm�b��ԯk[�橴�
�|�V'�M7��B��ي�91��iu�cK���t;�X�Tٸ���5��xRX�\��vC�������^�z�I��'^^�i:�w��]U�k����n��QzsYѣ��<Yh:s�T��21�X����);N��A*�PD�]U5(������uR��@U��䌊�߶��2;N��O~�c�.��*�<v�� ��{��^ս��j����'���kq�|���M����8j��\�~��|2'�wa����ӟ�,�GNg����]��B��$^��+�'�e��`�Gob�[�����+_� Qf$��*)� y� ���� ��h� Fpx�:�������on}�������WOѸW��:�y�BF8]e�N��<�먩�Ӵt�ɣh��\Z-O�Ku)2J�����8�~���{vf$盳��<('�1����L�����ѝP���|�s����&<#3N0�[�� 6�P��<~����Mg��?�?�eDm�I��ϡ�¦[�B�d�#����[sut��e�<��xS��3�%x�WJ�~,J�Kr0~Y*��T�6tgfn^��L752�&�L~{��5���]Q�m5�	���0�6�ma�����
��"L��,���%P6����nf̋�ox�c7tw��y6_ l���C(/�1��кLd��� 
0�c�&��C'%nb�qP�A��fX��ΓgG��bp2�l���.� �ٌc�Rowj�x�I���̄r��\�jU��#���� c�@��h	�Բ֨ߓI�����B�!d�Q�Н�-錬VjMyb��4!�c�MjYՁ	��cv�O[�]��ԓe�ʕ����D���yр�	�	��>�cȧ:�Ͳn,&�yDѬ~������Pq�0qF�ƥ��S%@_ǋ 7DM�~����@~�c��H��+	�:���m�5w`�KÏ$*�;�#�ą($/��L����lB���~�O�O2$U)Ei򫈰ck�Px�/��ٷ~<��d�C!c$��|���9ʴ��^t��7gy��;6ܿ��ଡ���Luib�2̞*�U;M��81����R}���c#�9f&,Ǒݿ�#����<�� ���Lf;y���ZT_?"��&�9���lV�jǒ�~�lO�2V�I�'��e<�s����-�*m��A'�O�1��c#��[����p,̀1YOǓ5�F��e�͙��/&#�,`�U��u�SG�u��g�D<����
� ��La*�Z��� �t��2CZ���x�y�yQ�Ճ0�aF�Q�{m��o�W�i����+��Dʒ7�wfc$G���9�3�r�Hn����yp�L��-&`�J��zc��m�*�Z��K�-)� -,��P��g#�FM��n���aţ��W̭-��H��&f���f4@�@B�b�� ��=�7K����1F�2ӓ���仗yq�|�MY�O����U��Ԁj)&/���9����&S(k��"*�Ь���
��j�#��0e�o���rcݚ�Q���9��RY��
0���ɹ-]�zc�+s�<���y�r\e�(p��K �O,�lI��E�J�D�g�U�r�gy�1�7ڃ� ����<w�X�:����j���c&v��Ƌ���ܔf8�lW�)��9b����H����#���Ĭ�r]��?�C��,�*r,�*\���FQ�n���O��80d;�v-�=�1�Io2P��,�,zyjh�G��0�l��Я%f�,aSgH�yl��f�J��W�/DRJ�>R܃>Ō9S�2��u��/�b�� dXq��Y�Y��1�Wħ�:��כ��eu���2�\��+1�-	,Pr��c���U�i[<��Wˌ(�ΒSO���č�b��d��0:�0��UP	>LJ��0{c��(����0)�|�0IU���/S:
Pm7���yԟ��n ���Lc��A������fԼ��Ŋ���t@�.	5� �I31���@�7U �vo-E<r�+�y4�P�3�UU� �F�R�̦[S-�休�tYr���0�>Ŕ��J�(���Le�Ų.��\3m>yR�9�|��F��x͔? ���}1���?6�l���UWK1�r^N�hc0o�IͶ	�A3���an���u�<wG+�شq���d� s�d���0R̐%�dB�c4/�^�4�c/�M���1e���%����y`�F��y1]�<Ց8ʖ;3�N��������{fR�����1��8Ʋ��Lʛxe��iR��D����&f��
���sY�'\j��L9�*L(QVD,�S�V27D�˹=��r���D��o���ӵ�6s+�!(�[�Reim�/ن��[�c�k-�j���)�<����Gǥ�&�t�}��:y�����;��y�V�@��ٿ�Zʎ��h\I^O���ϥ��[�W�/X�^�w�S�n��5qp�8�ڲOKϧ���UUŪR�yP��#�
}I��p�F}?U�0>����>�\]�'�l}�<}UHK���{c�-X� �tm�pn�/&���=���s[Y�������q(���<.��N��ޠ�N���6�^���u����c�gm:����t����2�����ȫ�c�gc#�JS�3>��t����m��h������pwT�t�V�S��g�D<���B�:z�S|�>���z'��ۺ���nV��ޑ�E�N˔��Z�J����1�g�� ����{���َ�i��[�O]�����.�ץ���Ϭ2��-+Y�]U��s0����ӑ�l5��%\	f,�t����KݒnN�n�[JՋS�l&�f�K����t�LFи�ו�c%�m� �O_vGJ����uwoT���!s��ռ��isHc��.�VE�+���"�����gM{N����zs��c���|p�Oh�	�C��;�����������2����<
kEa���N�Z�n���Cݻ�V����J֧z�<1G���ɑ�x��dD�]��,���m�8Զ����Σn�6m7JҩVan�]I�+�Uc	rw<��c�Y9��ߢ?�|N�������U�.F^7H���è�1/�����Ӵ��K���B��;�2Z����~0:>l˥�����x ��~/��Ir���x(�5px(�9��|u�:��'_�4m]�"'�a�^G�y`�HC�%]C�dVfRA�|v�_���_�'�������}�ױ��4]>�Y�u�2u�W5M3JG~��[�_U�5�JZ8�ˆn-Q�o���T��Y��ӽ��t[�c��v��qP׽VY �)����^�Ʋ�'���q����N��zv�R��#�3:؂i͓gN�!$��J�v:C:��V��"{��N����s��uۏj�]מ�{��}��]#��~�'B�:��a��b��է��4�n����x�����'�߄]۱�ۻ�Z���a���JŦX��)��5k���I����xV*�s��|]��%
{_M;�[��4�u�Ig�Q=�X�B�����������b���Y���{��ñ���G>�jXc!�,����i�L&��x�Q�T���~:v~��˧i{]�V���%�i��6X�H($�v��AJ��cS�� hj��J����4t�ƱM�r#NgO!���;T{�35h�1��^����v�[�?���jy]g�]����*x�9�6ve8���CZ�t\ĝ�5�+����.�wY�_�~84�u}��I�w>��a�BԾ�VG���%�'��I�|Rձ�ct9 t�~n��B�m�
�}��ObzZ�(��%��kU�hύ��̂d�6b��`ó=~�ݚ�i�}[�=�{G�{өWWӳ:2��}�>��]���j���Zn�cF��~�꜌�m;�)\��XvԱ�uս�b~���npk;��>F���|�'��A"*q�_#�fS؋���ڽG���٣�sE�� fmZ�=��������Q�����Xk�#v<��x�/�_��f=��X�E�'StWLwK]�#�w��p�����^�jT�ξ���ީ�1r�t�Jb�Z���1��S%e����������-˷��,~ЛE�44�G*�m>��'�������2��Y�����쾔i�^���锚������a�~�Y2���!G�M,��@c�;��o��������r�)�u7Pۧ:+��}:�Tn���&GT�?Uu�V��+�^#E�t�FY�)������~ �9E6MSS�����=
�E4�W�#(Aܧ�N���$��1�ʉ���2
u��^���RI?�b�@`��X�ú	� �������޷�xٺ��YR��2��aʹ��O���E�DAI��RvU�Kz�o�hM΢!���YT�� d����s�r@#U��YG�,8�I�r?O��.�'��C�ƶк���7&�pt�|xgb�|'#�l�̞R����n@Wi5d�O��j����+�������}�#���b���J���ܼ w�q����]��n�ձ��tfD���A}/S}3'V��,�P�4�t�P��9���"��y�#�ϧ������*�N~�#/�`���}��	f�I*����O!�z�ʗ!J�<�b��?����.������?�N��j���bW���.N7q���u���ݳ�MU����9Z��y�K͞����y�P�+����ە�=OF����5t�u�9��%'���+���"�Y���~��gZ����i����7iataA[�7{���7l�P>��g�n����O�������}��_fBK�h��=���:j�:��u4Վ?�W{d�OaSO���� +ĶQ�l=gW]뿵z� 3� ���CO ��=��pI�ژ� oq\�/��GZ�4	+��׌�'����'�!����
�Hb�c��������n�o������m�]c���:'7?��	��i4�����k������C�����9�4�j�|3t�7���e�{�wt�_ݿ��&���	b���jV��=ZUV'�hT����?���AS����������7���c��]�=��v�г4�-jPME��sͧwAs�����Ǳ��u�]w7�=��']u�Rw>����Ur0����Wӱr�ƣ�-ѭ��v�M���_藲i6�ÞV��9�H7�O�z��N�ô�үi�k�Թ��m�O�R�IYN���`e�mH���+�h1�iS�ۓD��S�!�F�����V��kPw��9��0��^�g��薷	��ئ�p�U���w������w��as�:�Gn:k�zZVֵ�̟ʾ_IZm��Y���ΆGS�d榣5�v�L�>MR����z��lt�T�zm�b֣vJ���LeK&:�M%��Wbe��*!���luo�N��Є���Ԧ�,q�Z:���ژ�~[P��=��Jգ����Βt���Kڏu5n��m��}��[i#�On���Ok3����M<t7T��T��{��	-��q���7'�{H�����R��7O:�B���̥�C�ڢ&��B�Uj��*ɣO#�KMa��rFDRvw���9�Z�追�On���ݻ�N壋N��%}9;ċ��O,��uZ($��W%7˥�U�ݵ�Dw��ԝ��]�S�	���F��n�΃����Z>��/�K�,���5l�ӺK������A���D��E�z��_�g��-��Wr���2t�ҷM)DT�mwK�0ڽ_��y��y�UuI�@�r�WR����wf�Сڰ܆]$I^齵�-����S�4��z�Y�Zm�M2`Z��19�^�������?C�h]g�7���{M�� �����.�'�x˦jO�Һ�r��ԺV�����H����W��j�%�F��_!�mZ��:���fշׇf1�ԫ�1�w�1�*A4�$�:���4��7?��y#l�ϊ��r��Z��֣���V���eTX�b�D�n�b��&9���!Q������@���ݯ��=����tev�^�;�֙؞���hF:2�/��lJa?��⨆D�g6��	�cHi��>F�0���m��z#���[k���i���-J�ٍ՛T�i�:=I�ԣ�����*�"˚�6��ԝѨ�n�kz��|�KF)-աX�NOٱB���E�fx�	;ㇼ#�y���=�{D��~���+��6��)�����β��5[���3���UӅ�ƅ��L�lg��F��r���$(=l&��>�|Cm��z�JqxSH�#R�/��ĕܩ��/�U>k��iY�9��U�^��M����[zOf�{��^�Vx��)?p�����J�U�V�#`^�����k����w��mS�z�#�G�m+V��;MԽ}����j�Ybj�j�)|�K<��9i�3��]m���A�7z�D��Т8|�q:V.Ġ�~��gPLvM�� I{�T�h�ڤƲ΋X�K���v.eP =(˅Вy͊��u?���_�'�N�tW�� d=��Gn;z�=C�c��Mj+�Hy�GY�ƃ���n�f��ٻ�E�_�]���ݚ��S�jF�I&�4��`/�gf�0!�2�I% Q�?s�WkI�-�hT��4�UO��1Fi�����?{+/j���.���a��{����:ov}�����|}�e'\�YC���;�a-"�21z��npp�V���uL�hd��|H���1�C�^�S`�v���4�Cl�����ܱ�C7�,�Zz�W�����\����������֩���6�ڡ%����o(�X�e�����#f�����؏s5�/��O:wC���g
Z�t�!�-S����cM���z����}Le�,|�#��'���xil��j�E����[�x����coX�M�Ze�=i���O?����ŗ��.i�A��RW~kj|yﭕ�!��-���5���:z� ��b|emBni�#��;~S�ag��>��a�Χ�)�{�t�j����h����z%k��zNl1���p�*�N�3�c��G�9��XX�v��[g��n6��2j۟^���+��ֆ�n�T�
�3J��;�P���',��L�v���|g�?7���v��fHki���b��O4��@���KI�UUo�Tw��}����gT���^�w�Q�f�����jt��dju���	p�\�c�]��-:73&�ϕ��KbJ�g��zEȀ6��ֻ���o^�+'�|�t��Pު����]��?a��e)�K?�o�-��v�\�lա�V����+��,�g�H<!k�U\�#��u�ouy}G�����{��߯Y�R�:O�z��zx��{�F�+f��u�Bah�����zX���(*�����z'�Z���C��oEޚ�ɲ�0W����`�s^Y��)=�GT2:{�)fP2��Q�ΕwfhW�޲���j�Z:�o疚,խ�1��$J�;���;��[���zֹ��o�:C��i�F���v��ֆ�����.n���'�(V�Ș.|����T��1�)7yh�o��li�����w~�Z�z�Hc�N���JЈ���	c�(yY�*6�����q_�~�v��h�RFY,۝�#�ݙ�IYRe�8�+ifq����{���v���	�z�Mh��/Wu�T�n��>�֐�mJ��V��k�6&n��ĳl��﷓`�6yoL��O��c�:l�n�2������*$� �dW�s$nJ�"+�{�!��6_M�J6]���+C���,��^6"̲#H�\����{J���ϸ_kP�o=s��������E�!��u�m@��@�Μʥb� �������Ӱ�G���ݚ��sPУtj��/��P/������"Q�,��IEj�a�U*�o��OtL��j�#�sW���o��O� M����~��5>�i:�z���u6V����j�=������|���^VF�)����x8m�3~����:�>W��ܪ���F`��8���ʪ�s��H���{�&�m����?�X��3E�2�䐬	���);�1��u[��?h�A��}��Ι����GV�����T/t���:��.�関�!�)����?2��h��Z����gg� �㻁��}ro����q����B�V(�!@ ��<�� 	�G��g�og~��w	�#��!����Y_�:�S�N������%� �uPG��|%��P�����h�nJƼ#�����$���>���.9���������>�4.�t'�7������.������ֺ�%l��l����i���\�0�7i����ƹ7�� o��g�ɨζ-�{�b����׻�0�����z�v�5���x�I�ir���8Q�O+�������{��t���N�wsR��.2��}��3���-S?2������mc!�����ΜW�]ӆD�=�%����قI��jE�+����� hHfCʑ���067*������V�*	紐O!����pT�]��^�=��O�G������-k�ښ�K�����'��|�:>��Z��WX�H�p>e�oC�����"{O��٧fG�������0Áb=���^�	�t[Z���Y�?c�=�-����(�����^Fps���:����3;��S�{c��m;����,лi�m*�+IFj��APfkz�2�\����x�����Vh����[�f?S��rÁ�.��˷-���?��@zU� �8�u,�|�FS8�n.������7��ٿ�V�Y V<����?�+	Y�����������^�,;L�k���pVke�����?����z����(,��y��������~��pX�1^?_a���c�u��.>��;5$ᕈY�^ne��?���M(�s)��_aH��O���-=`�"w��s���q�� �d,�h�P��n�uj|���<ز��}� '��G��̰����3�IE�1��9� ���g�]%�KCM꾫�a�����r�U������I�s`m�Q�ͬō6���ؒ�@���������*ci����s� /ow��?�˕s�MV�:NگF�jF.�~�C}%jꙉ������#/Oiѽ��r���<��d{sj��(�i�g���d�י�n�9�VfX� ��G'��#,�Ƶoh�IfqDOp��/<#Ui���3z�T�Y��'��oj^�;iۏz^˻]܎�����_K�}{Q��;o���V�n��=��?Bj9�_Qt~N~������5t��&\�e��}��@z{.���u���Fێ���G��&J��i�s"G���D����ݯ�N��疽z�q�oH�LMdh��+?oo���(fd�(������G���/���W���
{���'�fF���CK�� �n�������7���R�3���ꎧ�mp4����}SQ�=�\�l������� ,άk1���L�v�B�cK�?i_�q�jo�a5�ug�||��@�i�������5�W9ye~R�����N ��b��T���������}�'��{�����n����s���?O{��z���q�z��d�Ot��N�cbç}���*jر�SM��O�Ȏ>��&L�ٿN�o�NQ�;u�=*���c}I�y,W�� �H�b���sl��Ҽ�iS�Y%�D�E{�ۺ6������iZĉAK�Sku%	$���}v�j9�-HEv�!�~�C�;���~��9�^�:�������v��W����[����5(�O���Q���	ѷ��||�(�&�F|�|<�3�-�w¿M�^�F�M�=�14�\յ��Q�4ra�k��A��
�"�fhTv3Ƅ��~u�{�lC�7lZ���^���T4-M��W�g��=#�h���C�RʯǮ�B����OJ{i�}�{^�����\�������wk}����I�bjX����J_O�d����3���ffrK'k�����{#w�z>��mmf6�"������hc�S�<Z�̯��WX��?APyg��{�+�[v���%M[��@ex���\4Zu�V�U�YKY��sH�v&���o�����k�1a��f]a���ev߫z6=N5���m:�Ν����j�x��ssp�MC`e.6D24�e�n�i����O�:�����F��u����P�ܥn�&f��x�'���'˚��Ѻ��>�ٷSm�-W�Z��|����J�	��7�ev����4o�0֜� ��ߟR�yZOp�_E]n.�׺��+Нa��������JG#g;]$��7��z_��Bt��^�H,�{����;ww*(��^�}����ۜ��G⧬6�G�Y֣Ha��>`8����4#�hֱ�7�w{!���W����o�WW��4���z:��5��}WA^��ruM_Y���-��� ߎ���;fS')�
sO��#z�=�oE�g��i4�١R�KGO���� 6,��X��C �s��]�ۛnCoO�X_�(W�-�"���F{ �ҙ�=�8%%d�3ʎ���LgO�/d����ﾍ�No�~��}Ե]c����o~��[e��.6~D�MWOҰ)�;�>���9U���ț��|.��v��ϥ�I��]�Z�ȴ˺}َ�FD����$��u~|�B�PD�#�3◢�Gn��_p�$5wޣ.�OQ����y+�|S���BG#'�Z>8*ܗ�� V}������/��3c�j�m�?������s�fJ#����~�Q�z��E� �)�s�y���k4�_^�B9��9Yo��n�Q�����X���LG�ЈO�C?x$�9��e��{S�rt�� l��ѻ�����m���m�9��NjQ��A���lu]f +@Կ����ɦ6L��ul�<'@y����>�mۨi�����3A��{T�[��A�`5��;���}HR�:g�9����t��u4��k"y5K�,Qܵ�����g`Qy�\�(ᓙe�;�}��C����� ��{S�{E�����z���Aꝫ��u�<N�ɶ���u=f���[I�[�O����I��B� }m�Cn�6m`��h��d�(�"̊�S�	A�i�KDXƬ���T��?�~�����}GU�V���ec4�KgMD^+P�Op�y�9NҬ$��Ϟ��W�t�:oAW�4�7�m;G�޳�����-5��|L���*y��?���j];�2�kQ�Z}F�����$�ݿ���{�p维�y?|�F����NjZ���'��,ߒ4B����q�?b���=q�h� L��vw�>����Δ�;}�����^b�W�.k�_�L� T�5LG;�����˯d��qԡKj`��S��c��n�
���5:k����R/�x�	�*�K�G�N��S���l��Zܺ�s�܎僫L�����ߧ��B;�g:+���f`��5����w?�=w�ߎ���n��w�jڞ���t���ak�CM�����t�5�t4�uY�7Qǆ�X�ci��zd�~���T+��5'�o��8�8|�7,�Ah��ʽ��V_Sp�iw���{3i���Yy���*�c�C,����1���� (����� B�������������{�p�k�����3�?�/NiP�������# �����U�hWv1�*Y�� _�U��'</�>��|z2'�(*jo1_f�(�%��%�q�����k�;��Ľ���/���U���n=5m���\V����G\���=}�� ����_���i�uzf��Z�["����m#���5�,C��<� ��rHk�o@H���K0�1CUV�\s���0 ����`#�gg(���n�{��:u�ru�d�c�tΕ�+7FtL��Ӻ?�zgS��{q�H��A��er2�n%��"����A�^~��%�� mؖs�=e'��Y����?����*�
=���AZ|�Eu^'�/��� ������
HRw��ǿ��ϣ����Y�]�����Ғ�[�Y����O���M��!��Zl8)�(`T�Ҷh��Z��!y�XēH�H�y �I��.�y�9������nº��d�o"	�'H�8��IO$k+����w��9��\r�N\"�60L��MC���YX3�����23�i˞2tB�i�[�Yd�*Oď:��l<�� �UfM�b�Nc:��^U��Q<���M�!�^`P��c#��?㼃���O�4���
�S��
�êp��*��l��ϒ��G�Kqņ�#7�#2��2'ī��K�o!oȷ�Z��Xc�� ?p"����c�#��1���V�c�K5 o�<�;�f�+����X�Fk\c�)Tg#"�/����i3V��e��P�~e����Y��D�r�J-�\�*1 ە �	!����P�X�K�FA/�ߎ9��+[����8�n �r�'�����ˑ�gZ7�I]
���(2 6��ǐBn�
�ǆ�����
�P��ڤ����"��l�r�=iY�yVGwS�,��f8�V���I�rM� �fC�/�u���[-[yo'uߑݗs��!DU^O9ʵg(��n�p�*�ܼ�	��}�30,��^K7���cȇ� �"ye ���(��e��H����t3ܻE���+�� �]�V,��j3�n�`�����'��ݠ^t�U�`�(�R�`_�B(ı�"�K��93��Y�5]������zc1��)�a�����7�nBOtV�0g�_��p�vu��LaǍ����z��L��*6Ao/��F�0R�TIdrU�q|�QUԻ����L�l���e��'h�)�4d?�in�[�c��tV�J8;��]�)�w�L�ލyUc+@Ш��N�7����v�O&0�fY�Q*�"�Ra���� e��d-<k�T��mٹ�ٌw�x��"�Ek(�=8��q��\�2yX�?��	o����c%�� '��[cT�d�*ȔI�\�P R
20g��G�0[�ZfR?��*ő�QѶ*U��V!����| �1�LI�G��Ux?sHpm���~��9� �M^#uOLb�$�|V��V�H#4�����I�Ѓ�>+0~�6��K��[!!�$.�j�fk-#$�4b�>(h�D���ĳTK��I�[�<���	9��L1n'NA�r!S�|��S ��+�S%��P��弞�J�V�
4ʀ�F� ]G%,a�7�4�ʗ��l��9�W�<L��pA�K0;�6<�� �c���%�/��ȓ-n��,u��<��:��,`Zl$�H�ArǃT�(���k㣒wb�Ⴊ kS�j��S�c�eqT`�7�R��z/�p�M�P���Fӫѝr91O!���h� �U�+F�%�g(6`�Ui+*eyM��-@|���u��tW�TV��HMCn�H����U[�z�f�r�>%�U@Y����R��؟Lc�7 �F:7&���IQ�E�Ǚ������� zc%%+B`���S��T��]g��%�8�Xw��p�?¸bݜ��³V0Us�슔t.�ݲx�4�Wut��
�NI�eWDe�G�mI
�jJ�Y�{�����"��@OLaU��=�h�f0uia5fi�̫�2ṔA!v ��º�)���&���ޣ��gz��˸f$�G�1�S=�$�YΘT�UH0�#%���^py�[rq�HWjN�Ʀ֌f�UV�������zSq�>�� c���L�5w�l�
�f�-��|�U4g������Ռ������a�gW�'~4o%��=��^*�@�Vx��OT�X�G.?���)�E��o}��٬y9�>*z6�|f�3Y{���'Wþ8��|���!䥿&�j5���e+��'�sDث?�3�����9ak�Zf���l��\z
��9��(��-\�X�|u2���|���1������/KB���N;2��У�����<� C�
 ff�pf��jF�mg'R�Z�[�C�ʾ���t_��]!�9���<���=�?B�G�}���>���=�����?Q���yԴ�>��u����1e�Ql����h/�?ˣ&��#�o��G)�@��m�=c��;֧��H�����^8N�|�!���|�Ԝ ���v�%�];����з��N���Op,�)��VY+�5Ot����X���^�{0z���_��Q�q�a�=%��jz-k4����nZm��xn�J�yB���W�uյ��mön5Ϳjn�Wv���>+q7l��Pyh�Ub9(�'�n��-��6��7Ι���wѾ����� �t��w�ٻ}	��O�o��v��~����j�'u���c�v�S���:���k��֕��=c��ֺ�.��}0��1��KeFx�IyPM��}#Cݚm��ڞ�׷FMJ$�hj�`����Ci�fW���Vo}͚�Ҷ�S��{��KlO�@H-jZ%y����srZ���8%b�"@�#����W^���;߯~�]�tƝ��ڔ��������6-���ؽ#�t�Ξ<�ִ�z�Y+(FK�UJ�.4߂/�i7��]BmGUYl$�oA^��x��a˧uO�c	��5H�j�F:K� ����	�A��e�H#�VŨ#Q �DZJ�*]Gr��'w=�y˧�>��w�Iߍ�^�:G�u���ǡ�;w^��Ʒ��Zv��j�9�="�\��ǃżq���Z�ݦ�^�흻��u}�����u[����E�"��!��>iYX;��@�j�h��3�������oZ��z76�ͯf�kw%�^'�mɞ�TN��GUH��e.Y�mi����?�>��O��=/�{��]��z��U��jz��EХ�N�\������33�M�+.+Mh�TV+����G:ɷuN�4�v���[�\�rFgvSk1�)�ʈ��I�@��f[᳭�����S�Nޑ�kCP�B��A+�-eb�����@���*��E����G��K�wㇺ���G����kˏ�uwk�����~��d��	�S�5������1�D��?2q9��^�<��?���߻�P�;j�v♤��խx�� {/j#�40ܦ���>�^��o��[K�f��>��E�mV����$QC46\34o-i��?���~��{_߭����v�����L˧�[�:��.��܁�`��6nG!����C�>յ���0��3tY�CQܶ�McR��_��`�S�F�~ {�*( ܓ�������:�kN��uIfҩY�vKl�X�`1����X���ݘzrG��ԏ��z+�]��o��z���Mj����k�'\��U���6���t�Vzgq�9Mr�MA��e|���}����ֵ���-v��q�b-ON�VΟ��aXO�����׉�j��xP06}��k�n���/T6ōof��+ɧۧS�t�`p�M{��}�l����1�v�������olZ�.��xwS�Yo����{��}Vz�l�:w:���C�]'Q����\�L����i�̖Fk�m� q��]m���������Ե��Ӯ?� H�5�We�հc0�_3^x�X�W~ӯ]$��m�M�u��kvIn;5��o�$�0H�v�ȍ�`�'P��dB@���`��=��]S'C�&�N��11uv�||��j�D3���͏�|��.誄�x��6E�cB���+�*�x>�,
���x�x&�իH�pN}�T����x�X���� ~a}_Y�N�����>&���j4o鏡�'*��e0�qԙ�ZX�����[ѣ:�1�E{L񬝪ĢHUK绷����G<���V@i$��9=��A��� ���}���kA�\�N���}��YԳ:?�Ω�`�X�Qԓ�s,��aN���eV�'ybFaN���6��Y��X֮%u�eW�K�aø����2���ʰKfm7T��E0;�4�VrJX%c$�H���3�O����웼�౻i��un�.���oE{w�ֳ!�.��Mb��H�w��l4����'��)��d��rc���]b��Ǒo��sU��xt�C��_�[р���,�ubSQG>iʛ #rق��雊v�#ZP	A��vW�&�����p�ݕ*��,���W:�'���#��Z����{�\n��.���l{��9=��4��b��x��>����=���jOM�Ι����q�����u ؝L�ۣnKӝ�����J|�,֖==>h0� m�jf��F>I�8�&���Dl�����V��Cw>�*���<�'RMjJ���0�SK���;BH
��bl��}���Y���d����]�N���z���wn���u�#�q��К��}R�m��#�g���k��(j�ǥڙ��jZ6��uMc|i�Pi�pա��{T������\��~[�|ʣ��a�x�����E�ڎ��t�v��������,i�+�Z�n�>[Q��ĺ���ѓMB�7�y�x�x}����:67D���;}����������{=Խ��=������=G��-��3j����d�/�>���6��Z"��/W�����nj�u]mَܲ2�fHTX[n�d[1�{�$I�;�c���ѝ/lЩ�j^��+RX����GXEC`��R>�A%N�f�w��F�����YǠ=���=�q�&p4>�n���Ԛ�_j����B��u0{�:�4�Jz�D�'�Zw-Qd�^��tk~t�]����]��=_I���Z���2If9#�~��ȑ`�H�i�F�I�D�˶i�R�Q`�[/�Ewf�OR[�ӣ�֣$!�O��t�Y%d�c�#·�ʌ���گ�.�{��|}K��WԽ��L�q���۶?ou^�ԫ���6��N���wcu9��9�H��&Q�����OB��FΒ�&��WP�E���K�kS�i�9"�3UrŤg^Frt��Z֘�z���k(b1ŬЛN}�Z?U7�䴭�ģ��b�QXӱVy]��x^�t.��Z����i}���t>gj5=W<�V��ü/C���A���?�>�mG�q���k����S//N�������� Y��V7����&]�&�6��m�"��Y�-���1MF5K�MZXa�4rD�7_��y�L�s��n�O�Ы��SQӡ/X��L� x̺l��^jv{�y�a/	!�{A���N��
�/�����ӝ�����_�}��:oR���V�>�����.����5��� E���E��9uơ˗��S�?K���ὶ�T:��E�C��T��Ln�C%YV�j�yZF���[����Ԏ����O�[3h�IݨEZ��5�v5��H�H�|ԎbyaD�����۞���oԟ�;q�����oj��v3��<�����W�o��/�1ϧ�]S�:�&��x��}C�������˖9�6��η|>n]gOޛR�����#�.U���Ҟ�_�z|�G%��3��
�a���;�q�{��[��m��黓aO��m�wkȐ��
kW��|��7ŚJA�Rgv����`;��Ǥ��wc�{�:kَ��E������t�{������N����r���:d�]W&X�IӃ3A��O���� u�m[�G�/[��N�m�ŧ���Ѥd�Yh��J������?uh�S�5{�$�H�9G�F��G��f��� e��/�G�5@u���̶a���d[�U�x��٭i �G���wy}�{V�Ww��~���y��{�����@euWZtN7m��g�a�=����F��|lSS*2|�6>N|��� ν�)ݝ:�*o��
:6��RWէZ�yCE�h����#�{V�E�(��el����u5jt� oڻ��>�Ug�Đ���J�<��Eg)�8���?���_�m3�����sڟG�?S�a�f��u*j�zv�2�58un���g/�-OI|El�u�}����JB}'J�dX��l��Ui��Gk-f��'#��p\R}Dg�^��V���֚��_��ٮ��	,y�i�~@A��=�N����٧au�b~�o�{�������@�v�Tӫ�^�8���G��t^��l1ݭN�Hb���UuL��Z�2�#�݁�~2hK���&�ܴ�hlI3<U��+"R��Ė����Ũ�i��4bU�YD���ѽ~uH(Ձw����bj�[ė�Ȉ���+/��"C4W+��U"��w�ou�½�ks�~�����^������op�B?�tj-$��zc�r5�;ɯ/�ǻd쯔��j.�G֩�]þ7dsh�mfi�'�YZ�#���֯J�/Ù�F�"9p�'Ǵ[ժ��nI�=��������E̦͙�(��Z(�{-�2�O�����Q�����m{�ֽ3����Et�]��:_[�@�N�iZ���ck+][&�C��)ԫ[����ԯ����ة�i���?��7Mƹ
�#��}C��R�)`xa�Hb2�ӟ�}V�Y7=�SS��j�"�jOR
s;�4�v�o�!̈c*x�QH��Oo�W�Ok�������G�?v8��vˬ5�靫�gRҬ�ݾ�������8��֩��d6������c�{6�����[|Q�mf�R�]��}?ʒ4(���X1J��z��ig�O��EkH�~�)�nɼ���W#[�uj��W�ZT��,M�Rj2�fq<�����P�A�Y�{K�52;�G^�24)uGu��[��]d]I���|�/)���Tq3�"�<MwK� ��ji7c�-�W�t��O$/fy�>{
IjR���Y|��<|v�9i�����t��K5�\��@,��?I�Yd�V�������_�����Ͻ�{Y��{��A��w#V�/�Y��vOCv�1��+�}P�U���Qc`_Q:�2m(ͤeK�fZnD"k��s�R��'�KG��+|�QrK5`��4�#��D��H�~����m��϶�;�W����_"��U���#�Y�H��e�V^#UU�y������z�}��"vϮ:�P��֏�9:,�����t�|,=C���� ����~�M O/Vck3��#����>�����ܗ>~%Z8*3:S���!���������;B����ClS��ߠ(�3��kvW�KbS��Rp������9f<A��ޯcK�������x�]��?��v� U�OFj�1��beO�qpc�꼣��.������V������ٓx�����b��;�F�V*���4K�2���s�F��)v���,��y#nVX�������r�,���{�F �+�/���G?_��s7�ޭ��i���ބ��ch]fǶ<ܟ\iX6��Y̺kI�_�y~f~��ս5=F;J�&�Z)�;�|�x#�����x�s�o�<ps�'�c��xC*$"�G��E��}��H�1��ܗu��ն�.�u����b/J\�\n��	*�N��1:oAJ39�2(�de�')��c�������?��?��?��]V!�q�O���q��C:/����N��{{��7��=�����^���]P�����2ftIt?MS��鬀Y[ԕ��q�����5�bH��n�4�5$����?��g��b�/3�9�������>�խ��Gvק�c�����k^��s�����yz��-[��`qt�ή�4�뮽��(5r��~�h�h%#B���&W��C<�Y��
�wz
A�G�x��f{R���4M⍏��;ye���X}M��Rsq�	�{��oi;��x����g�ž��`������a��ֽ/��˩4l,�|�Ro���9Y)}�Żq�Hd+2Ӗ?�7qGn�V?�ו��Z���C�����G��c��'���r�琒��G��������%�3�=e���:�;�׶&[��^��� cuu|�mo;�]3�ƒꞭ��5J������H\�}�փ�^�y���A>ݲ:��p}v�'� 9��RgU�J��>�� |�*V>}P ~�W��V�����=U���ԽU�d�#]�N��su�{ṲA9�����e�䪁��MR\QB+J�)y|��{#����\���㏽Tr��ݱx�~��}� ��x�+��麦3�j���ÿ'!P� Ԟ���������_�vz27��>��~޾���럱׊�%��s���� @��!�����<��e���W������l@�o�-�^ǅ�<�x�~��������P�]Sנy� _��̍�ϧs4˵4Lģ]�;d*q�	�
�"l��}��r>��li7c�2��� p�y�� ������R��P��O!���o��=6��hR�\�B����2Դ�\i��jy6%�����KgX����*?�A﹂>���}^������WTi��J��ڥ�� '�}� �3+KK6N���3��}?��l��H���#���܆;?�n}yW�P�6!��icM7>�䛽y� 9q��8����·򐵊�����Z>����<����Fz^���uIu�u�O�K�H������UҸy�GN�:ϖ�~�ս����f�:sխ��L���M���Ώ����ium�+�F��M�̝�ZI@֎�Q�ᾘш��9���#�f�1i���t�3x�����=�����~�@ 3�>�=�{U�D��}K��׽��+����������<�[��ht�'W�קt.�gi�\mD�Z^�����l���:l�F\4�Y�zY��t��4y$��w��="��u�L+cP���}�Յ��(��wyY>��6�W]릵�׶����d���]fiD2���f�6%d�G��ƥ�IX�z=�f�C����؏s}��������^���f����W�4��w�;s�CK�n}�m)Nv�����c��ҳ+�b�?۟PԨn���6��ݷn��N"�?�Ow�WQ�����5Y�d��n���yөս��7�ۖ�4�jջ��~���:�)"��^�4w��{'Q��.���Y��to�/m�����Q�Gw+���r%����N���C��t�q}=n���|=K�F�l}#^16��jt��y�?#w�z�P����ߐ��?U�N�պ,�g�:�mi��X�ey�i���M]`Ŵ.��>��{�џX��ۥ����w��u�h���-�kjA;Y�`~��O����Ǿ��^����{C��ϵ��[����E��v��xt���κK�cu�s��:�W�V����}Mo�}=n:���~�j��-�kO��]��WOԬ7��Hb{�kqج�xhB��M*��I�u3H�/)�i{�� W��}mbB��ؚ�XBA�$u�S�KY����kʱ��`F�9Q��� ���x���������uf6��>�:ǸZ�Wk����w9t�m{_ҳ5�B��]R�ɻ�y�ZpȎd�,Kj�r�CKzթjtb�4�H��+A�$G�qE�UC/����p`����v��<۱Ӓ�"]Fe�yd�U����ܲ��Zy�Mڇ�@FY�������.��?:��/ݵ�����_q�������]oT�i걮$��ȟ�ze���p���wz���������z��v'������ʲD�P�#Ce��	�a���2XGS9w��'�z���mv��ۻ���j*5S"����S�K �4+�#xQ##�u�/���b}�v���n����j�X�Z�;�==�v����tg�N� m[f�#3�oZ�`�cd�+���t��`�%��P�=(�i�X(Av�%��^P��qF�/,i������>!������h�).�Q	�.�nґ��ie~X<��H�nb�� ̚�������uG�m{����>�鮯�;[�����l^��F��kO�s�p�l����%�ZZ^u���4^a���Q���j˹����a��E~.��e�!���@8!�ި�|D���\_�2M�H�����]&H?gS��}CJ�r9��py�O]����'�?��}t���^�ư�߻�ѭ׽3����:�N�C/?#Wѥ��{a���7F���y�����t�mlϊ-�sV�^؆��Ҭ-I�F�]�@b�XeA��*��D�Q�2,jݣ��a�;���wЩӭl����f��t�X���W�Q�;$lȮ����dfr�٬�����_ԏ��a}�{��.^'e���05���?H�N��g������ech�-�S+S����l��gl�u�0��]g�{C��>�{��;Z8�&�FF�b^�VVtY$���(��b�K��T�������f���c�:���]�,Ԅ
���(����y�X�Vy+:����s���/d��r��tG��Z����e�zw��k:������rt�.�5>���N��%�l�[$���-5=cs�\JJ�|P�� ����Wկۖ]9����K5oLC���@�?��İ�P�@
�v'h�_þõ���m�Td�V�Q�V�Gi[����.�2�y<8����9�������P�������j�r�;�z�ci�~����Z�~K�5	����G��%��>8�n�?����մ>�h��h�0Қ�ڌ]�+-œ��O�Ux��q/�� ������ dޑ��i����5��Cm4�L5l��2�D+�e$2CFbc�B��%e￿�;�ھ����7�c�I�n�����^/M���_Pi���fv������լ�$�]�mJt�hl-_�zs�h���)Zz#3Nl�󼎝�v�j2w� 	��Л�y��GE�:���X�2]�.�f�E�t��$P,hݑ�0fFd������׿Ν�9��A�Wfzw���잁��9�Ұ��Ꞡ�Q��;+?�c�x�r���^6k�ׅ8g� R��g7��ĭkQ�����Ka���ջ��n[���a�O����X�)_�V?K�MO�;WbӃH��b`�JakQ�]Bx�0���$�����y?:=��Lz���s�{��ݶ��uOx�����J��4,5�ҚRt�>&n�7�N���Ǯ`Y�V���0��t?����z������g2,q���1��O'��04�"�;��!��9��D	�X ��	���?q@�Y�=�췷_{���ݖ�};�=���������0:��2�����r��41ރVĦN��fԿ|�:�څ}{N�^
�]�3�Y�	�#YG!�y��^��2p�|�kN�+��ʶ�_�쳢�Gy�3�%�Ǣ�y����ϰ~�7m{��w~��k������&���v���s�Z��Y��֝m���Z��i0�l��bFɍ#RE��Uզ��#�j��H��̟y
�������*~D�J�Q�#}-?��a�,#}
@�¹�O�9���Ykz�Tuf��uQ뚎f��k��u�]cYճ*o��ꚞ[�s�if%ތ[q�� �-#4�{�����8 ��g�!W�@UQ�{��� _�盢s�ܐ��M����� ��m���}|�~� o�����׿��&O�񡫨��/'4_����A���؏_J�G�~?�ϖǳ�����g҇� C��=����S���?�u^��ݨ�:���ؚ���`��6��L��I���dݱi�&`�Dz2�l�����n��;wh/�i���"U1�5t�� �9� w)g�,�z(I�4[����ר����[vC�5�V�Uo5���{S�&XmU��u�8x9,�H?�;7��=Q������:�K��9/,LܼZN6SW�f�q��8M噂]N�}�x�=J�_�۫I�|t6�v��&�$���:N���s��d���cx�U1GF>2���׫���cN�<b�p�ElB�̉6����Q��;F�MVP�^T�úe�;,'�*c�#�7U�ڑ��k��9ێ�ŏ���B$�Hd�)�h���du%YYOYXe A�ΥC4V"��yVx'Utt`���IVGRYI�H ��j�6J$�k�,�C!J$Zk��/�����vۇ�zdf�F� ld��(������Pf��{P$��2]�J��,�I���#B*�3�(\��JC�%�*�#fc#Q'F�'�c&��h�%��JD�h8��^-������K�S�*&<~g�v�#��|�������Sd����6�@��	�r�4�cU<ه&��%Cn�a�9(
�l�4��p�K�/�ĳ���Z1��6�ϫ�P��(�4Y����K�6��D-�1�/1�%�-f�[�+�1Y�8�FPP��į�y6^\'�~CVx�El�f��	$�]K�%� x/ �2G�1��έwUc�m'��%Ыl�]*7�Ř�,���`���j�"d\R+M��l`��2Ʉf �6�G6ܟLc�(�[*m%�)�<�x��_��6�tٷ�(c$�S���UKZu��iF�$����ظ,̠�%}1�.�o��?FR���
z�B�C�h�\��F�b ,d*�:�
?U4���|H��]�c��Tj�;3��u��,c���h�2�Y��|a�0?�Ǧ3�yBW'�hWy�x�$�)kAE�Y<�%7%\8m�
mtDi�V��RI��@,W�ަ�yq��b�6�HV0�(�f"�Y_w"ng7l������H�P�~;	c)oN
��ƥ�j��@l��`��:X�)�.�P�b%��ڨ�0�/6�B�@։K��E���;�~@o�=1���YO��۔x��;��+O�J�}
�X�`ԗ���y��r$av�@�K,��;�@U�PC~�]�1��|j�a^g\�l�o��M+?#3'#�H��YԀ���c��"�fZd��+-.� �cy!�~�I$�ըA�1��ScZ@�-F�dz�dQi��*o�;�B� ̝Ԇ2�(%ZlH�񷋎<L�(����<���ն��.�t������s��e{�%�y0G�~�v,a���NuHΎQ��eF#�CN �d��, �V2�Պ��յg)�2��RJNV ���TV;�ܱ���d8��E(�ܝ���á��t/2 �Q2��)�E�OPQr�ԅ,Q�MP���se ��b���c�e��s�5	�P���yU(��@ �FD
̻�0>��Q�i��@���(4fu_6��?3��	e �1y-���/�le<�jS� ��[
V�?�(�ۖޘ�6cz��Q�g���`�E�ϓݎ����Q6� �2%��Q�q�M\5[�UW?�����	���n����*�6Q����G�L�'#�\ə���ŏ�1U�r\}hA�pIڕ*Yh�B��!���e�]�匕�R�"3��,sZ���e�����l�зC1��̈��p�(�U��9:N�E8e/b�p�eddGˌ�&��_3K�9�Iy:N���'5��A����E)��[���%ݸ��nC#�\�%޴�<Af0��$*�D�9,���|��̈�� �G����Lb<�`ĺTD�S��n8���A�S�b�X1���[�r�|a)�q�rf���u@#��G��Ա��0L��ep8�Ƨ F_���)�y=��J�� ��rx�c��M���f�S��4F?�!��'Rͺ�e��1�|�%2��,2U�dD�JQ�`�Y6�c&�;��g��3�7n��N99)4�)�U��V����T;�ʡ�n�w4���h/t��麖~$��pս�e��܍[�l?�N��[6� ���7]�}1�k���KL��h�)���#aNr��^���N2�Lf�Y�8��0��\zc4W�zG��Mrq��<y�&�=<O&@�ᩚy�[(]��
�;���>�u�t�a����uV����(�S+��f�8��-KN��4�ZN���,��p�;j��:%��dp�9T|s���4d� bUe����n��n�6M'p�j�\�pC��p%�d+5y�?L��H>��zϤ?���T���������G�umB����c�m��Y�wc|�KWDzU_cAH켧P���˿ �v�N�׭�wes�ao�ס�1l��v�w>�t$ �6OO��g_�~����d_�}��dd�*�R��$C�Q�C8��N��kz�Y�u<���M�����GO�xQ�6Ǭ��mguMgV��r���N�f��B7� P��tf)�O�q�2/pb9U(�WGrY�q��ĿM�Oԉ�n�Z���7�NDFf�<��eYcvBRH� ������Y鎿���K�{���N��]����֏E�/J��,�th}S���c��TϞ�lmK��J�ʸ�˞��Z~6:K�� 5_\�>�a-��b�?#,�|�V�-Q��sFC�f)��&@�Wt��}��t�z.��ݍ*ӱ~=6� ������k0��9#�Q��д6CB���}��Ht��� ێ�k��^_���k�3����j�]{+�4�A3��W�u�N-\��]+*y�ՄD�t����=�?�>�h ��5$�t�hV�6$�:�5s�<�ZيK��^أ� �q��v�o[>'v>�R橷�ø-m�iEz(��7�0�Cd�F�F���bV,�n}��P�z=���V������.��=iԊ[SҺ3��3����jS32�������ʶ��	-�mz�ԭ+�;]�n��/��:��m��<��Q���,��Tw�^�t�U�R���8�t�{/�2-:�~��Fi$�a�9
Y���+g{��W���6z�E얃�(���Eze��U�]/�z۹~�����=[�}��0����JZm���𭅑��aS���|Un�ϫۥ��ڃ�CI��\�V��^Ē5�5w=�B��O��� �q�Q�6N�ͯ��h��n����Z�"�+9�Yx%X1�"�0eQ� {���������t:/?��Hj#ۮ��5����ס{��� �]+��^����O��_;$N퇛X�γB�>M�����v�[�m}=��Y-(Af*�'VF ��=�7������<t*|�7�ԃ���1�K�\@x���p �{����:��ΰ���g������5zӫ�=�t�>����t�i���Y�޲�m?��!�a��ɒ�q_�����#����V���m��lEZ����sM�8�5[��ȃJV'_"�Hw
P�n��}��k�e-���ݽ�X}&D���՞�k�Ud�a!�>�]	^��#�Vv�?NctoGt�_��p��Ϋ��G�6��'s{��x��=K����6R�]����"Y�1��YX����I�p�3�|�_	76�V�ϧoui�եԻ�:d��d�Bk�X ��Q2-�\�����%_�m��;�j��(�R��5�~۪�Ru������`�����ޮ�u$���}c�=��<=G����e�w���i���Sk<'�W8d�;G]G[��`NQȖh����GQ�P%�mױ;֧N�y�[���(�����{i�O���e��WzR�3$Q�;3Zw�a�E�d՚����Wy^A��pp{��OgX��魢kZ�w:���=Y�kR�[�}���y�_l�
?.�޻q��IN'�:�^��r�jB��ln��85n��M2��á,��}p�����h�l;�����:�F�n��K�I.��I>dx�� '@ؿ�vg$���?찒{Q������Y֍%��l>��~�������މ���#�=�v� �����7�q����g��{;���ڦw�7ҭ]K�i,kYUng\Q�-N�V�>���̼���S�M+P�ν͵E�f��?��EӞV_	�v{ǭ�j�tޭQ�x�^CF�[�i�ue���u,~:l[T�1"�u�E��'�{��4N��K�~���[�1s_�?r:w7O_h�K�C:f�۾��FYbv������5�Yg�.���叕�I��km��5�W��b�}ѢN�]f�מ6�T�`�5�=�6�����/�cl�ݺ�����ݺ)C�j�٠��UE�\Ң��3���i�`0V�X���9t���O���6���u�ږz�j���ܾ��޺��5��t:��1�yu��2����bc�jk<I&W�M4G����=aGJ����;��4����Y��]�"Z�>T,�(N������-s��V�#��>�E%���i2�%Id��ePO��GefO�^�}��u���o��Q��_��Wj�Mս���Og��ߵ���ug:f�������7Sb`�	���m����m��ö:��~���m��X^���G�N���I�Wp[��f�?�V�,� {$��Ē��g%����}��jz6����.�-\�[Bg�H�j���(�ZE2�v�B�\�U��,FO,�8~��z3�wz{��=��z�����]K��ݮ�� ����S�o��8�����N1�Yt��uON�N�o��Z�!�Ke$%�c�w�[�9Ck�����7�t���[�w]��%��Y{�S�Vf���jEfh_ʱ�dn��#`�:-z].�Q�FH��u��[[�>n��<CC�R�f����#�Ȓƪeq�;C�Op����Dw��o���Q�n_M��ԺG��_T�N���s�'#AN�a��S.���WR��� !uJdLd�b���g�7�kqk�B^�n6JF��إ,%G�DccɎi����/�GћӼ����KnO_M���햗�%jP�y��y,$���$��|Mk0�I�k�7�y��{��r�?Q�� i���l}�z�z6�n��MJӴ�SV����pe�z��Ek�����ɗ�8vi�_�B�J:/Ӿ�|@��Pt
�-Yt�}sLYlM4Q��r�X(��(�/���3F�Us:[]C��M����c�6�4P�{��C�V(&mF��H-<�����@�<�s��k^�zK�׺���O�vZ�������OZ�s�N�����n��֑�퓽�z�a�u$�a��z��-������^$ϔ+Ԏ���M5���ޣ��lRAv���hkU֋�z�,J�i�b_P�%x^8�����V���=ߢo]Snǰ���A�.h�~r&��B꿓J��q�R�5+��9�o|���g��Τ�p� U��[d�?�z�;�ۮ�?��O�B��'N��������e��3[&9I�tSe|$|Ek�VΏ���ZRK��Ҹ�F�2�3�sN����G��"�7Cp�\t�l�:^������Ӧ�F��a*�f����,�L��Y�����?f^�=��g�>�{�л[�^��}F�:�!�K��l�b}[ֽ���2��J�ɵ��[R�����z��ͺ��>�����4�f�}Ƿ��Sڸ���b����)X* ��֌��k� ?�Nnun���uŤj�T)���	fy̩n�4�'�J�H��$]�� vO@{;��������K�#�{��}hu��S�Ƣ��h{�)��ZwS�|{U���Ng_L������������Ǟ,���Uҵ-W��S�'؛�6���I��U�����<�
Έ���d����8�{�J�z������t�o=�*����A-k6U�V�����f�[q"B�����>�=�k����Iݟp}���{��i�e�gv�p:�J�FQ�}%;c�+ǣ������<��["��-Z��o������]�h�Ŭޖ������I��Z��j�R�	��Z��&x�#]���D؛N��P��F8�MB/,��
Y�Վh����;��G��>+�������J�f���_�e=/�}��������#L����3�|];Ӹ՝�%j��]�f���{"m��o�ro����sԂ?��XڴT�y>�V�U���������į�f�n���V��#D�����ՙ�Ov獂S��UQ�^B���_�eӡ� M��FT;��zݗ������'S�{�,}#���~>��� �F���?v4ӕ	*j��ꌃĺ�Riо26�����;oB�CVY�ݧ_Q�$V���D�%��F<�X	=�[���ֵ�{��T��n+�qi��/\�V��,l$�M9���"06�Bk1ٞc�FO��p}O��W�������qt���;�헫e�v��z�M��t��_+)m�]_U��z�&��aJg���ISk�������N�o� �V;Ҳ�V��V4���N�6�H���>^¢H�,����/�-��-�&��6�0�RI۩�HX/̱+����K��w��)037�晤����E�O��l=&=�{;���i=K��c�.�Mk]��4?����|�/�Z��el����e��JS#���}�����6�hn}�r��v�N�]bo�&{R(g�!�_�b��	/Ȃ��� �|bj����"�o혧�P���!{S8yR�QU��q�{�k�<�gi@��]��}��M��\;��=���#��w���=�:;��*j���ݨlXޘMSB���ɥf�.��Kb��
��'����so�t�cj�Hd�A&[6P��$�fh��4!�ǁl�	17 ��m� ���턂��f�醟�ҕ���BQ�,qG�d~X��^Nάû8���{��G����W�� ѴL���X�:~��:P�@T�#��q��æ3ej����rrJHk�MV��Tɨ��bF�ʎ�@�I=�/w�'�Ӥ�w ?�[-+W�H��aȉ���GЊd��=�����joo�Ů��֓�Zn����t.�tDtWw�E���?��?�:O�1umC�s����KF_���S3+VWXcc��_Yմi�����dc)���rÇ�vR�0a�B�?Iq����qp�'�e^9_��UJ)��G#Ȥ7?������?Tn��zv]��_^u��8zi:� }��J�^�u�,�z�OL���;e�|[<���^�ϛr�V���Ů5!R�GH�չR��FH���ߖ<q�"��^H��v�f�-�������w#��_E��q;��l�U�:� Zu�W�?��.��jZ泗fjي��Xʢ��ȳ�!9�#*�%z
ig�I<��?�I?��s���>ߠ� �� �} �;ا��a����kў�}��b`k:7b��u��v_'8㾉�uޡ)����K�Ň=9e;��o�������f삽�{U���?�Ó��Dz��7��&���2����O���d��uΣ�'�����uQ���ZGSegOU�4Դ�|��Z��t���yzK3񥆫��*�?K��}>�ҬUDjO�� I�x��ē���9�]}��S\����[|�O r@`���/=�Ӑ~�[�}�{o��˳2�'���W��C�5�jj����fi��Rpjet~�ڹd�]u^N?����yb�Y�eݱR�k��w��Q���C��^�V<r���^T��'��
����J�^�M$�yIe��
��� RhX����~�G����?���`0z�������֣�9�n����a���#��K��1�g@�Z�c��O..���3�3ߕ=S�-��|X64	�� � ���~8���r�kA�h�{���<��?�G��~�����>�����|q���Ê�+��r8�����%�G�����9�_��W��#,`�����p�Ѫ�+}?&.�Oj@���
�o�	gC� K�����bݯ����������Y�j8 ������ׯ���$4�x��	��#fƪs3.fb�j�3�6 '/�w2V�p��d��ǮH�����sGX�I�j~�����������?mC��C�M�8̕q����Nũ��;o��/���g���$'<p=�����z����8�����?o_����6��\7��ꮉ��I]0HedQ��e�99 �� T���������I��p���}�$/�/\p	#��]�i����H�G���?���[|X]-�<k����9������t�Ԟ��.��Y��զ�~�����y�%�5)�X�v��7'����8�w���ߓj+.�JU����ȝ�rD�n��@���;�۾��'f{���}��G7J�������~�S����m��=�3_�WM�l<Z,ee�J����Y��� z���]�sx�RR���*Ԗx����H�2 � :�q(��#y��4*6��?@�����n�pY���c��h�<B[��b�֮��;{i�|u6'����=��k��^��L}[�N��*����占��轾���ΦNɍ��.:��N�E��F4�օ�Cs��s�z~� �C��Q�-���]�c:�&�f���ef�y6 c
��S�E��^���k7����ܭZ�{ԕ�r���F�$Hdr��l�os��]E�1n��h짺|�v�^�=�9x��;��������罺�4������S���Wty��NNF~7Pt�7��VE�l�SГbT�.�[�fE=�?C�q-OyIa�޺���N~]�ѵX�H�b���({im&��U�7M�Lk��*V��W�`��+�kL~�e"_���J�,P��Y���=��}֝]�\�A�/e]1�zz{���t4������M��Og�	�ؓ��_Q�ZzV��<�7i��z��i���o�ޡCC�ԍ��mpL���4��ک"�l�Z�<ҭH�c�dră��^5�-�.�%�wB�Z-��n�Z���K�T��dQ�������J�������ބ���}C߾�����`���_�;;؝7A�=�{���X��t��w]�x|����Ii���4���Lk�<���� ����n�f��7��ҡ�z6���'�w���QI
�V����jSb��$�8˳5.��֡����[4�}�� ����[��k��j��R��`Q�"��GH{a�m]��?Կ�w�9�]c��]?�]��gM��R^��-?U�4=rX�x�״��|k[%Vm�[���3�
��ӿ���1-~���l��4��0���4تa�U]�Yk��KRv�e�H���hd�c�oSz!��W˾v]�:N���%����i'��l���8�h��X$@��%Ic�8���+�p��q�����G�_D��ƞMt~�aiZ�y�k.	��/��#Pg��v�.�v�<���ٳ]�4:/����}X4o8�� �i���8�{j��}Ɖ��7��8z�H:=��3�Ff�v<\p�Xy�{�8������޽�a�_�����j����~���]���#N��'V���t�6n���5:x�3MҰ�%,�����A|J��%��_Nv~��̴Q��)�۵����ok�(�-$�i��d~��zƣzo(�vnzAe�*V�W��U�I8�UE��)��;�0�o�'�w}/�}��3a��j�齺t��O���k�5��*��5Lkb�Ӳ���Ym<�L�Dӌq��=s|^;7�]ݶ�?Z�-F�Pڎ��/<W	�
�S���{^7�'4����jG�6�u����:m�.̦��w��n�e�6p�v��^T��o�9XzΩ�� lY�3�^�꽜ǏVa�Ji�w�l|��o3d�q����2����7��޵��K¥,w)���{���<�8RG�$��_��v�&�Ku�v��������~R�r�HEW�~�f�v+A��l��S��tR{�����
tnlc�c�D�Η���L��zj��z^YY�L�hi�8���k�O�EՍO�Nm��Zm��t����%5)nԗf����F�Z>�l/i-�h���_�?Ҿ"�E��ȃZ�z��鏟"Ju�^a�Uz��P��I!�%���Ϻ����R:˹~޺W�n�~������Hw��z�������5<'B�5�{�qp僯�GQ���n.c��0șY��I�1��wY���5�д�Q��k�l��H�,��9G-�f!�;)�߄���пy�i���Ej�T��W���$�Ѕ��I�nx{�riƫ�����oUui�w���A�R��A՝�]S�z��sR��<�.F�<�ś���r޴rH��(>z7���3t͵�+��xnF������^��ʄ�~0��U�[�]]ٺ������C�ڞ�6��4���<%����)��0��7���`�o��j>��{���o��^{p�<mG���랡���9�O�uޥ� a�����T���*�ba,z�����X3�R־��ڝ;�&��jP޳r}.7���똑+��I:�I9��� ���φ�oY�濹��u5-Z��`�� �WM�a�-8��q7l���T��@��w��(�� p�.��w\�c��ѽ�����ѝ��ǲZ���X��.���t���ύ�g�G�� i�6Vy'Nzy��nZͪ���m�V��u+���x�g2.���AT��Wp�֕��hP��L�ݥ[��{��;$`ݏ�'��)�u���^�u���zc�}��6��>�̦��Ӻ��m]���4��իi����P��3��ݳw�s�����F�RX�<���{X���#`DĞC:7��
r�uZO�m�H��}@v� �����{���9�]��E�^���������6�����[�k8�G��x���lXd��?Ve���д=6u��ċ����~�@��pnYd1I�D��L��:���G�;�3
�>��*�������̓ﻲ9�`}�TQ��'U{��D�K���צ�ݺ�^�-�՝C����yI�\���Vxat�ZlMM���A�<�d���&I%-�'�O`G���`z�����>�v�EQK�?����_\���&�Qf>��w�G�}v���o��>{x�� ���L���?��s���-�_�b̠$|$�w?����zp=�?���>8�~G��2�WTG;ɓo�||�I'�|� ��o���?9�9$�0P*�~@g;,��Y�o���7;����~w���o��{�s�o� ���H��G�S����nʦ���#���k��{��-�2ճ�Ô-5`����v��?eݦo�Rѕ�	;,I4b$�#�@}�����H�!��,�kZ%���_Ӽ-OV&��L��,(|�/�:+v7
�+w�~��F�K�)���k�j�-��?���Y�6���N���h�X�'mBI�㜥
y4��f�z]��N�^�W�n�ʦ�r��1��[�qC0 ������{Yy���ΩR�X�(��B�h��әG=�Y�d�� �G|rOŀ�1�6ц_;S<���i��\�i�֍�i�ٙ	�N�Y[�J����Ԩi�m�:q	m�;��b�hf��� 8�ܑ��}�l�K�uMc�ۥ��t)j*SVN�A5�]�^�I?��j<Q��d��2�R*ƞ9d"mM�-�ŋ������K6/ F�`�L�VF��ҕkg	 VEw�Y��X�qcV����S��lȑ��n�hdO������oLe���g2�N���a� u,� ߳8����92��uP:��Bː�|-��ψy���9�Ɉ��$�r[�`�7R�u��΢��+�+�*���m��A�0�J~Kک�$��TqY�QX��+�r��e �Ic*hIfSD�ޜ_���o�ATA�~d�ܰ��Lc*�g�<jLxUr*�z5��2�r��� �;� ��c�1y(�=��4ߊ�lv&�*�~�
��W��M�P�d&0W�@P'/+$ %A�/�Z��-o"'�Sd�Uu�$��,��P6�Ō<��Y��I)bi0��$�O�@bT�!�Ϧ1��DZ��R>Eɡh�eE� /̗U 0,hኞ@��'����oQ��*љ(���p�}� �m��1�UP�C�VaE�~(�v�5f"h�S��J����C���!� ��T(�� (l�B��m�?�>��f�+8ȰD���d�q��(Ĳ(�	;��� )$��y8TPN�J�0Q&:�]�,�m��̫ *���7n*�9
���q>D�q�I��P�i)ra1Ƥ�0]���2W��Ae�)��Y	�^>7ǂ�)*8js,�̥���Gt+?E�>i5C�7[ng�.܁6 1�W@bc�JC������G�b���X�K�Y>��SU��I�t�o�GiI%8އ�[xބ� ͈R�1���U�Y���*�^F&D��͛b�X�O'}�1�vYը+�i=<lQ�k�@��
% �'�曞Jȍ����#�S���%ky\(�M� ��*�vO�ecG��-�iEI��>|h�&�w�>F+W+��I�.�r,c���mYN�D��P���F�76 rB]��c(5s�<a$��Ȝ'�f�Jի�O%h���
��߸~C� ��x�VW
���,�:Odf ��<��!�k���S&	E�����5vyN���Ķ��w�g�³�o�5lx�BE��|)��*��r"�G;�y���D+@�Q��9���8� �%����H>Ė݌{K"�q�Ƽ&��Y����Ƴ<_ÎU��(�6�.��d{>E�tD�`����j�'�%Mn�Q�� g3�j��*U2��{����!�@9l6�?���*�Va�q�i��?)�ԇx������tP�����3�6��
�;U�D8�f9HI\�T���r�2b��qST/��X;+e�Fǂ�Yx�Vn!�Z�X�X�� ��-FF�����>�#b��T��A�غ�c"lVx�J���T��%W������m>M�NL�`�\?��e&�r�s��[!d|l�i�����p̜ATW%���*Ќc��|��-_�D���@{���� ��~X�L0)Eg(�d�:����R�j)G27 |Q���>�fc9y���Z�ޥ�������)�}<� 1�����O(x���o!%��TV��w6��$3錎ˌSM1�Vz��/ǘ	AQu���+�n�v +��c%�r�y��ő�+5)���PlT�*�7w�[f2$�@1�8�x��_�i^E�� ����6�Ǥ��!)�5�;Q�
=1��tE�A��(��ee(v݌���Mb�V���!$�F����`��FRL�0T'f.ZͷV3X;�ؼ-X�FP�3��B���$�?�	f�Pi�ϟ�%���xc9]�� ixK���OOʍp��E�����UY�fȀ�D��b&�/M���{~ֺC36�8�/,�>`�'�W���6CƳ�.�`�vfc5��z�d3�pӉ�Lٝ�`6-7'�����}�~?O�s���'x�!M
��.��z�edt���d��QVB� �]i�}-(]J��!Z��fP�/��n-��i�c]÷G���`C�?%`� '�B�%r����7�=ڝIiuX�k�����O�Y�H)�B���vyGeP��zQ�\>�=� v+�i��������б[��Bk�?�Ը<���N�.��ѹ7< C�0��_�W�����$�t�[�@��~���ߨ����XA-IW�z8(.�]�'L����N���ƞ(�-#iZ��q�7!���Z����%<��!���~�����W��|�t�i����mS�z�N���6l��c�k�NXt��r4�Ï��cP�z���F�"��ӡ���ci�O=y#��j�Щf�>FI"��YYy\�wS��Mr�z{WT����"�� '<�Z�v&+$w�dD�;�x��9x	$'������C��Y�縧�7n�t�:{�5]G#?_��h�8�ɴ�
e�W���f��2��|\�ۦzV���ϝ�k��Č��ZxR�U>���A�vw�3߂��O��aԶ����A��=:��:�%��#��W�sG�!{�}�rk����߿`��w��?�>�u���w���l.��ZΡ�=����cf������mV��24�G?
+�0�þ9�v��%��W]�cF�5�N��uh�5�sy�e�ej3�#���,?�KC��nښ����m�z���,L)��5�a�^Ux�eep���%W�2���{���g�s���HѿL~�w�F���F�x�u�j��12���e� ����8�&1��a�H��A���ĄSٗ4Yt?P�S2�ѡ���� �Ɗ�wrKM��0 �kS�&�!�n�}9����� �2d�S��I	�#�}K��K~���T�gt���cݾ���M7��TjڇS��ugs雃�}����7�S��
b��
F}� �Ș��|8�c_�{�a퇱�[D�WS�-�:�t��g�bGt��!�UKv���1#>@_]T�����[�����ҥ��-��Kwpl!�I�f���v$d�>Ot�f���&��w#�:u��i��z#�OG��z���d$r05����Xv�;W����T��z��C�i8���cu�o�v�>��3U����f3.�QՈxt��W�߈�hW`�{��y�N
�B�M�+ԞQ��H�ǨL���[���2���kK]�r`�"ai=~�����A����:'ۧht�+Q��ugC�T���]?�� J�u�sU����L](�%����M��V˃�Y��)t��t�1�[�����X1-���[��<q$j�'{����t
d�Ƽ�Mkwu&V�_�O�:7���%]L�,�I�&C�'}�2�ڝ´���Ϸ�k}g���7V��=S^Ӵ>����t\��Y5��<^����t��d�3��>Lk�U'�uL|�d���MOco������sקf}j$�Z&�u䒉ק&�9��� �4�O�[.<��>�ۻe�M��$��$Q���4v��L����JA*�Z+�����l�O]}��O��ct��}�{|�΃���=Sڮ��@�� r�3���WS�������7��4��<o�|�r�sr�n���m�� Q��s|\��3�}�^�G�.�^Ĳ}p��펤u���u�c�����Δ잔� SiYږ��-gj���X+:�kBx��Գ��,��g�����e0��������{c랼��n�����������#7��粹i���ݪ����\�t�#�� �MC�=+=c:m�_����u;H�Zv�ӭM�Juc�N��؆}7Z�!/�]���a��Ifw�!3�3(<����ke����5X�o���)�g���p����V���V6��y�g���=��)���n�ﷴ���{�Y�f�S��E�|��л+���X����.����O:�%��U�=��@�?*6�˺5^����{�Ɵ�ޛZ9�T�)��U�WҢru(a;Y����N���[���hu�D�ю��&J���k�� .��Ԕ,�5�qȊiRJA̽�g`=�c���A����a�=���;�ڞ��-3����=���ҩ����OQd��֪�c4G#'5��^�:��S�N����Vꞛ�5;�uK���%o�Դx+Ή̳�")�<uVֆ��xa�>OZz5o�˴��;�en�i�_Qi_��~X�/t�`H�Z!���x�dg�ꝛ���o`�9�i��E?P���=3����3�X8:�e�N���t��<�Y�:�Z}��7����O4da��f���ݩ�[?r��S)Kcn��Uը|�2>�^H�j�i���M�̪��4.��3h���V����sK��CB�ձ�X3X�t�I����j��+4+�$sv2x��:� �����������c�m���\�loy���rj]����p�����h�-lvv�-��ː<X����Q6�K�B�"궟�6���i�7%F�8��u9����'j@����enF�űw����uk�V��v�����:Tk3v��MSK�U��	QȳV13�@�B��w����������n�����V���j��e��ן�~�{������L=g������ſP��zfD;ϟ�O���/�_������7pn�ѵ�Wէ�͝-�J��a8���TN�->4�(y򒤑���b����'H6f������`���;��c$�Y0���u���3,���X�ڡ�]ǯ�_�߿��}�{��N�w�-ӽ��g�����������c�7�3�A��bj1�������8�8`b�ܜ��&O�ބu��f����N��t=�z�^�$d�*ո�XZY{D�dV�c��I��Ω��w�#�^�jZ&���9�n=WqQ�A(�̶���N���,k���3�&(�|�O��7�/�������������������eԽ}�}���f%a�ѽI������GtN����Q4X���A趁�-��o��f���h��mm�H��K�R?wq��R6���y�lN����S@�.ܧ��`CKR�:Ɯ�v��P<���mJ#`�h#R��/�å4��Ǭ}�j���N�莜�uVr�I�=A�����n��кI���7���1i�#Q��>^T^"��.������ۃA����k1�Jԥ��Lu�-�)C�`Ր����P��PT��ݽ#�%9+ˮ�ZkܙRx�j4����"²���E��(k�p&��� Mn�������B���W����7B����ƋmK��m�)�N�X�pz�^���R�t�=?*�/NƬ�w�V<u�����O���F�!�����O�I٤�/�0NĒ:����̫�^�������im�
�J��)$�#�X�hp<*��9��2<�yp�#e��}������=a�]/ߟo}����\����3�:��ӝh��_'6ZFO2���*�]�2Ő�4*��x�\z]�4�]ͳ��zH�TЭ@��0��:Z�X^ʲ��� Cޑ�s�e�t/��k^�-mM�R�����I�(�f��f/<sT�Z�c�O�W^�4m�T�gJ�;�n;9�?i��Mu�F��ܜ�Թ��Һ�O��æ�|,M5�\��uޠ;����Ҵz�>k�b� L�730���������Mo]�v�"��k0�5�DKB�F�)"�d̬�M�F�3D�$�eWJ+i���[{O�N�U�mG�4�ZOdW�O�<�	��U���/����9}�?O/�o�=���Nw��|���P��s�:2����޾���~�N���\:�		I](k��lv�1�O���Q���Ϭӹ�Y���=AW�9H�P\�%�E�cT ���r���d����{O�L�Q�k��םG�/%���݈"��'Ҩ\���C����׾�=�{��onx��5n����7O��j}��z�S9�v��v�^�&���yx�x#m`Ŧ\� ���������{3Lкq��	7��p�Jr�)ʳVA�[	,,�*�f����B4���8�>7n��5ޥk{���6�ũ*Ԯl�k�n���v8fCS��)[�<��4��}s�~�w�}�uv'@ewQ�I�Z����z�:P�,:g��V���/�隆F�rNp�4�ޘ�l�-"z�Ԏ�n���ҧ��K��j� ,��J�	,�4V�Ҫ �eHE)<���>�^��}}Qv�&-gW(�g��~s$)�������˷|����O�n��?z�U���Σ�n?Gi�f�����t���]��k���}E��T�|�ˮ*BU�mF�.�w�Rc�UЭ,u<� �Ѻ�2�$E�r!�=Ï��2���9̲j�y����td?K ̌;OԜ�ܩ�ە<f������А~�uv����t����v�,gdw�0�Z>n�������t�G��E�a04-'%7��Ja�%�O�0<��^���$~;}�y�**Gf"��H#�G
��>N>�0<��J������=��3�&���V�7M�N��jڧFv��4������g%�MSG�U���yvr���y���BY��K\5�Ջ�Z��(�z����� ��.<�1�Yi?,�Ͽ���9�ÒO�ҍ_)��j��97�k� j�|1�nw;��s��?�}��3絮�w�=�sڮ����,=3^�����V��Pҳ��y�&T���Ī�2dL�'X��\t���eU`�+�����*���o���G�P�Eb(�P�,
�##nYH �O��J��ϰ>�uN����v���\,�'���t��	��2F�}g;]�Ӳ�zGP�̼2�� ?E�%��NX�U�����g:>�޻���������ݒ�+�;{"�]����=8�AEq϶���2�K���xO�u.~��}�tw���=�k^�3:�A��^�����2zf������l�7������c�� J�O� h�l�y)��u�1HoTU5�ѦGr��!+,�Y����Mf�����³��+$��;ƥ��+")1���S�"������tVY��{:����z����V���+��IhX��tWEhb����N@�t�pW�l2��jfd���b��3/�x��^I�|�y%�݋O��|�a����������?� �1^���S�"b63��l��X$ϔ15���$�yn6עێ�"N�S��s��q��񟂻�#���ۖ��?��~p��-q�I>^.B�aι��y���E�rA`yw ���F�b!�R^C��)���|��,�ȯ"��}'����s� ?��_���?��e�,�SȊ���"�:UJ��!��G��ћ� "�5=U
�L������x�}s����Z�W��+����?�����=� Mt� ���q둪�v�L�JX��|?���zrL�Ð%�l|��{�t�qٹ82���@�V�k� ���sϬ�J��Md퍔�v< ������$����h�D����i]5&V[�:wSL�w6��)���<�݆ɹ��H����{UijT��Yf�h�QI�v����s�>��蚮��bO���"'�c���������3�k� i4W?�:[�ǌ&N���Ӧ)��#'��.p�R�ۍY�	!�U�GO�[�V�[L��RغI�d�_+'�!Q�3�UG�׬�m���=��m�5O�<s/b�	�%�>�_����?����M;{��ڎ�ugI���n��t-���m�+v��G�]O��\�����K����rrq���u\�f�lV��t���2���m�ھ������ �(ZZm&
l��yd��8�.��W(�4W���C����m��KB�X����Ԗ��rq�A�YbH����	�9����e�}wӺ�/r��=����{oӗ���i=ӗD{�즕�+[M�{��f�P�P��^�MK��N5���?� +��ɸ[p��'q���������7*��{C�d����.��~���C�7@w-,P�pi��i{�4��n�~���z�B�P�����t�ooW���7l}�������쿸�u�>ܴ\^��_]�K���׺n�OK֨�}���^��ֺV�����z����}+�������`.Q�.��5�~�������B��_���o{n߂n��m'Z5��8oGCP�"��l�W̳o�� PҴ�[sZٓn�_m���2���Vt��58�D�c���g�RW^�w%sv�/������v��ѽ�j]%�?�ˣ��w�ν�x��տ���G[����"�w�j9��,���|��]=24�e���t*���̻�]�X�J}~�V���X�O�u�5�҈�!vX�ң�'gwd��o�7R��F��v�[K���_Uy�Y�'� -
�$�l�b_")��N�;�ڧ���h���o������I�dv��}���'H{P톤�����i�s� ���s��4��m[#Q�l ���tX�.���Α�,����鬶%��Ϭړ[� ^��ޖ��Oc�8�>"F%c�?[��{_״���mGS)=ѺV�*W��ʱ�q�� �w����goy�;���j�^��p����k���-6W���~��'Pv˸Gn�hJ:U4N�Ӱ|ٽ4��,h��:Ja��+�1k9_t|)���������w`�:��.��d�B�n#Y$�;$�/kLd[0�F����ԯ�{�v%ڕ���5Y�,�߽k2��r��HP��X���%Q��]�>�.��+�M�l�!��� ꢝ��=�z��=k�i��?պ�P�.��Z�|�=ޑW�ȴ���V̶7��Z�u.��]n���v�0�Z�f���<��!��)��G8��������4�Pm����Y�Jfu����D*�f8�ʢ6�pM*9�:��O�_�5Ol���� ���I�/Nw�]9��b�gDuK�P����G霌|w�vgǊ�/�Z�T�H\����暬:���V�#+W]6[PDcb�G5�3�0�DTUo�N�|m�CnAx��:�Y@�b]I�ٛ�}2C:W��"�7*G��q����-�����O�?���];��.�`��ϑ�������ؚ��`Qe��,��<UĤhڍ��q2��`��t��oB�/�����~V;�� ,@ӿ�l���W ��Ԡ��S�b���F����~��Zl[Vk[gQ�φ+��ڧfߛ���O�G<O��J#��U{w���u�>��ٗ���{*�p�i�t?\�n�'�:��Az}��'��ԯƵ�Uq��H��;��K໦=��o�f���۵�����%j1��4�l؎"���b�*y#0=w��]e�tm��á��a(��;���rQƷ�5��´�'���X��t���{��}����]��wt4��g�:��]WB�F�կ
�n�>�Ӱ��{���)�q����7�P��ǧQ�ݗ4����>Z�����ԝ Y$	Űe��)ݽǱwO`�l-Cj��_nѿ^~���N{Fi�2���� ʥ#U*=�+�6E�7��^�{��=��V��q���u'���i��}3]_^�2��굅r#ˍ������T�x y�Tl�H�f�����U�v��u(�j��

��^�Y��C�;�3���]ymh�.���g�s�����-ȩ�:T�5�o;#��y$�Q㈅t�e��݋�ٟ�w|����;�:�}��\���;%�Y��2�Q��� R��3�j�Ft�i��8�qf�e��̛o�s�.�]���	I�6���'��X�X*���A�F�U�pǈKW�����5mfh�tL�h��K�H.�&�h����E����TsО��O�_�ߣ�k�o���� v{�����}{��5�zJ�����N��i�� ���ɞ1�U�D��ˡ�a�]O���ޫ�!�z��*l]᫧��:��R)���#_$�VV-�pYTo�L>:U��m�u�I�W]N��nhĲIV$P�7=�@'���+�����M����G�������a�ò���H��-1�4Ε���MKQʛ�|�}G:뙏�)`	2gRj�ɻz��4-+N�;�mj�Iz�ؗ�Q�D�y�@��^F�{�C}�D��+ljw�=j��o΋�׉#fC��R5#ƌÇ�DiF`� 9y�/k}o��i�� d���3��:�wF���W+S�5'TMjZ�o{����kK�a�L�:��
=��XZnsA�Ԓ��ebĸhч�5����g�S�93&jf��t�СN�����Hd� y�O�L����^��m���q�5�uL/Ժobpum;�������\����t�i�6ٙ�Y�5}^e��Tq�>�^��VGh�H��*��'z�B�����υҠ�`�o���!��P��@y���ʏd�'4����~u�}W�uU��Y[�z?C�pzC�4�q��0/jֹT��2��d�Y���u�(�O�ǲ��%�����;~Y�ôzʵ�G�� � ~TzTRO
>���:������ ������c� ��������g��<���G񍳯$ 줖�����?��_L@�����p2�#������S���� ?^]����<��~[�9����'������� ����>�����?�� �����wo�@F�w<G����?��z������?��a��|�� �ԝg��1�Xt�S�����!|���]?N�!���=CS��uNV#�hyQ���6�c5W�f�u~��ܺ^���i�迡_��D{	�K���ꧾX��Xp9�?�HߛN���;Cxϵ���CUk�	�S9�$5kh�3�#���,��9*3�㴞�4N�h�oW^Q�tu05W�:�d��k�L�+[[�z;�#�U��>�W��5L����>X�=�����f։I���0�!��B%����a�ݒ��.�(�Q��Eww��{�we?pjin��s�߻��JN�g�B�S45(�b�^��1$C:�ԙ�.��^�$4��>���$\X�����ǌ�b&�L|&
�o��A����{Y����6&���=�<��%��p%v'�I�7>��;5�*p���ѫZ�Ѩ�a0 ����2� �}��z�+Bg���H�"�$(o�2��O� qRX�gX�\=��e�+�"�LeJ(r��Q��H���0kŨ��tg,I�n�ɕڜےL�x�}0#v_��-�T��Y�@3+��	�g2�^~\��	5f�|��cC���o;b��9�c@�*xf��<t<��KPdؒ���KR���%u�x�+��8��r�-��+[6˹]�Xƻ�(`�ש��%g�	0�F¡j�Cn�@<�ȫ�oLc�L���B���-�(�@��%���+v(~��Lb���*�p�N̖�wFS���ɢܨK|&�w#v1�E)/*(le��"7�	Z��.��B <y�X�� l��P����Z��\BU7E�������wc+t���JʢQ��\#l H,̡������L`d
Lx��7[��vZ;q)�H�%wN���X�R+AH��)�<!X��/�#��u�܈,ؐ}1��L�<�N(b�PR3b?s�W�y�>7,��O�1��
�gyD8$��)���4Ve�e�F#b��1��gvqy���9ed�ى?`1���?��Lf=��+��q͚aT���$ڏ͏6NL����`߹�}�RL�d�,;MZ��K��U�}Y�ERwm�2�vZ�ԏ0u�C:���h�R�:.Μ�o=�?	�Z��4؄-O%�^1C՝��EM����y1�厈����`�T�U���Q����Q��رc��Uڤe<�2�ѣǉ��E 4����'��C9b��5�1�&�T��K�G ��v�:��yq}1�~rw��%��.1,Ѩ�Ƈ�4+30� Wr�c͌
�U�zJ��_5g@Z��~Z�_���Yɫq�U�;F<j�5rXU���`Y(rdI�NS��(��$�� K����gS�M�yy�<�!<B�&Fr���QU�x��c�h�|z��������?�-�&��c��D��{�:��PH�Vr�(�O+�Q�#a�U�V��J-��m?�cv�[���]���'=�g����0�K��h�ֳ��2I����'$2���*��zch��	%�N�U��䛗�ZW����c!l=<hh�ھN4��r����$#>��Ռ{-U��*��J�ԥ��r�ގ�,�@�1��7���tN7�^�Iʓj�ە�$�lΤ*�ן�n�����.+l�?��&�ɹ�+}�:�p�Ta�i��+�y��	��iv�7ݪ1]v,N� <���G����5�Wĭ)��Y鲬���'���A;�A,a���$��r*Q�wGs
��`B	%<�rݹ0�e�o�[��@&�<t0�n;(v@RH�����[�+6Mݣ�f��l�bҟ9�$�+����1��f��I)'!�L�@����Eؤ�K}7���+���TG"3Dt8�Z
"�sl�{4�pNLG��#�&1�Ah�g)z���@2&�hh��.�D r%@�3MĬV�+���kHL}e�����p�8�?�%@aT4cB�e<��*��Tx���j���m�A���v2>�D|z��4ꕣ�&����.�|Y�r�LaB�mGNK6Z�M��7U`Wy��EQ=���c!��j�1M��#;QX+����J4�0��c�r ���gWD�)�Y�%��ɣ���0�B�T*���Lb@��e�2Y*��:F�C��٩��1,X���?�zc|{���^�������^II�-�3� ��ޘ�Q�}��y�,)d�r"�5��Qi�1��ᘭ<u����<�Zgb�i7v}��V��#�K��1�����P��2��,�l��K�f�g����g{��G3:S�);�X�|��|+�-qqc@��s	�d-E�*��n�c9��}��&��LTk��ʬ���� C�qB�8���f��a��:�J�l]�u�G@�]'*y:v��f�����x�:T^)�rG�0B��[�jZ��z���]�N�*7tsB�9� &_|�)�Xz`G���t�?X�kK�hũi�����e�T?ux�?��ʟjA��e����z���.��[T��w3I]����u�Op��:&N*���H@c��:����R+�9$�T�7㛵���vj�������� ����w_Fo���:��^W�n�rbGo�N�2���eG��_�>�Z�t����srr4��h���=+�1V9��.FGL�e�d�O�
9yHq�xR{n�j�4{Xb]sjjf)���p(��^Aާ�w2s����ѝ'K���jf]��MZPkGʓ2�*�^�m�n��Ъcv��=��O|�B�n���E�:*X��.�u?Qb��q��4Ύ�Ͷ��%�[K�ى�� � H��o�BI���,�I��ߴ�S�^���ߎ;�� t�o+CTs)]�&���)#ߺďI{��f�6�@s"�ֲ��/;8t^I����>�WG�Տ�H�i�m�;ä�Kգ���e���鸏`|nZ�w��ތ����=EkP�n�5yf�!�j�Mq��=�Y���8VP[�^��� �I���.-r��C�Y��瀉pW�=�D~��y�[݇ꭁ��9���<���jغ��ޮ��i]Q�N��-,.���E0���Φ�5g��5jY�FƘQ��P�=;�_�Mx,�}ab����--j�E'�޹�On	�4$J YZT�N�u�(k�ɥ��У:��mX�b�o-ԩ�z�$GHl4�g��Q$��2:G�΍��i�g��Zu�@�����Jh:M��~��u��<z�:���~���?V�_͉��o���յ-�g7���k���2�*K��G�SȢn�)�-s���3D<�t�ݲ<c�3׃���}n�M� �}^�MU�_��ͬk�VB,
b`� IOm�V�|1��8��k������}��M�zK���{d�m=[��ޥ��y�q��1�֝uӺT��w���ruީɎn�g���b��]\վ(��;��x�]K��P��WuJU�r	&�[�R�$IWNYbyd�@ϛk��=u���M�Ө��ϖ��jY�~@[V 	-�WdORZ�LS�%bH`+��� �z;����/����� ^�d�Ƽm�:��Yg@��125�#��� 
�����"q�}PU������Iu�3Os��M^B�������2	�������u� r"5lB	����A<{�~�9�ߎ���ߧG��OQ���������]O�^�us��V7%닁��g�:>mSwlK�%�.�q����|�<|Fy5�+H��.ᤊg�S�)��\;K���g�}$rI<��[{���j�wt��eY�������Ow��I�JY�9\rxe�B�Cm'���=��[�NwC�wO�������՛V}c]����7X��5̗�^���zw/1i�X�~e^U���Mq���G��[�zn�iN�a�v���K4q�Ө��1�LL�#�)�D��Ò_��'\ꎥ6����-G�$�K(��q�[�I�d�^1�X�wd��{U���~��ޑ��KJ�Ū;���7��%��n��:Y��J���uy��R�.*.���VLm�V����-׾�}j��Z��S�g�J�L����Vn�x ��W���ξo��t6���ڕy5!	����%�"�O��q~�@���`Ԟ�������wy}��vw�}��M�z�#K�Q���� ���}3"J����w;GV���x��j���굦�1a�,i�Ofv��j�<�;�����Z��o�#Nջ��:l�CY����b(����<m1���{��ޡn���liz�Ҹl/�
��lir�(-����V�;FoO� bz����~���;����:s��Y�i�a�j:��ӽq��%�ݯ��-��Q��i:�Q��sK��Ŏ�	�.��ǽLqk8����m��kni�'R��0ި�]��
�9�M>�fn��a��j��#H��1t2�E�{>�ݶ�M3\ԮlMfyt�M%��й��K�eP�U ׎�
P7a�v&a���뭢{�鮴���h�=�N�Z��Y�]��~�7n1��34��������l���7"yc�-?)yy�Ӯ_�xjn6�f) [++Ԓ���CB"%��!XbK$2"21��Ck��<Q	^9L<E:܉�`F%������gxyV(w:���x?ߍC�^ܻ3ӝ����l�;��۫�1:������&g�.�dv�&k��t��їRa	��K#P�%LCn���X�e���o��ŭ����ҵ���X�a+eH.DK9Y<���FH$��~�hX��U��2�OUҵ�T�����[R�y?f�ݱ�b�H���{�������=��z#���솭��n��^�;ف\�険��������lt�]/36��Fe���7��E�S��ͬj�tlCt�ߚ}�*��w�n�G4o��4�	<I2F�In1�_��cW��f��6��������Fv��a��+K��4�B����$u��1e*���/�'���^�{��n� vk��m�W�rz�?K�^�w�:S?�}*��� ��X� �r�3֯����o���>~b��z�Lz���ը"�S��9�I�߭jhc�'����cW��xXF�,�������FU�^��^�R�5��R����
^���a;�{�I�?�!O�|2F] �O�s�=��};!Ѿ�������� c�Q�����	�z~��t�[ur:n�u��K��>�����c֙-��c3V���=���� ��͎�
p黒Z!4�)�1����� c=k3Q^�DA�!{s��Z�ԍ���ZK�t�>�Jx��M�4_-J[s/��1�����Fn����O�z�:����O{h����������=_B�o�����SS͟s:D;�ڽC>x�Z���:r������x�iZ%-[i�}�kv�j	�.��C-}N�؍�_�z�����1U�Q���%����k�Ɨ�w�GG��$�Y������"L���+�'���*w��H@#�W��~����Yݬ>����L_l���.�D������/N�� �lG�_k��Oԣ����l�#7'O�+���w����s�[�z�~��Z���d�rV�BKZt��"�"�	!O,bxah��n%�q�{�fl]�WM��*(�K�g�k�2��)�g��v���n�Z%*y܎��N�=�{�?`�#�T�oٽ'FԻIݜ�]�����#�d��H��+�:r��Y���� Q��������t_��i���^�/ٺ�7;�/ZW��øJ�H\C�Q²�����[��|A��N-_�J��qu
�Q)*�b!�
2�	�E�J9�B�ew�z���������쯺~��.��ۣ����W�����.~=��=��;�})��B�Ů&ޖ�ϵ�ȹι��mj�u��P��;j/*۩c�f�-rl��f�U�	�9�T"r��������ֽj�P(�Tjr���P��+�*b�z̤�IQ�pK;��������ݯT�O7^�P��R�.�:KL�G�e�M;Q��q1��S���$1��J6..�0��	�6�Z-�,��� "H������!�ߏ]��$���w�^��֔a�R3������p� Y��<e���=��5ݎ��f���1z�u��u_j���FN��5*�']�.��4�O��OKn���N��sp�49O0 �V���45�RY%��;3�T<���}q9�Ȍ9k�ާbX��Q���Ы�ʪ�G�#Ҹ���$�{��#��P�M�=�N��I`R]�Mi�i��Y�6�;k��.�w?됸ֳ�=7L�#D��r���{��m�eD���ye�2�|F�u!y�$є�WڲD�c�� r����O���Ϡ��>��5=s���W�mWZ�:�Y�/��j�A�fk:Y��+U���Kj� ��6P�]��P$W�+{>�}��� �����e����~������~ ��H�~?�� ����}*���|�?�~ك�X����~G�� '�;� ��� ǪG�g�� �d����]���E����)���DK?��|� �W8��9����?���['�^}� �ٿI��>���Ȅb�]9֗�«�W�������;�,�z�1g1}��k�Ls�L|{�>�ҁ�x�?�`{��4L���,�nb'�����3�iX���n�ӭ3 Ұb��kR1�ǒ*�u���6Y.�3U�� V[VZ��H�Ǵrē�@�Ϡ ���2�Z+�!P �$�,I<�>��I��������\3Z^e�KUi����e����m��}y����� 9������#�_��h'Q�Dx'�������� |v���C�<�N�e|�x[8z(m���r�m��/� �+\�Fz�HG?I����ۏy���$��������2Q��j�Ro�̝1��T���y��p������~�
��lZh����� ����g������� \�q�-wJ�ዥtm�qu�E���2X�����X9��
�'U4�\��6����ޱ���%)?����� ���'�=rV��O��w �	�������#Oӵ$�װ%6L��i�MR�d����N.3�WB)�{�߈�ՓQ������MȂ��1�[�� ���?�澍�4�%=^����?Gia��x����O�=�h��ۉ״^��w���[jZoL�[u�L�zEtz�����]r�6&fh��<��]�\W�-/�jtK�{�R��t��~�M���~Z^��∰X�G ��B���>u��lݩ��p��;���K��=��_�{9�ƽ�8��3��ٿM=����w�r=�����#��IԽۀ�=�{��͞ov����N��=%W3Q���r)�V���H�]�R�U:��)6.��u	7�6W�OL�]KP�m)"[R���+�qr+�� �L�G�w����ڷ���ȭ�m8�-���:s� �M�*�=wIK���Ƚ6���=��C�u���ݎ_s�#�v����f��O�.��>��.n?�� �}��~��3��j��]����f�$�B�{��u)�O�]����V7���e�k�=*n*)�X&:ތ���t �5�'����%dnnz�o�;�-gr�5h���u��^u�C�*I�#�+�Ѯ��KS"��α^VUT�>���{��Ό��C��P>����s���7��vZ}�����eiZn���ud14��4n���j�c�	�4�CIa�A��5u��CV��>ѣ�������55��V��8d�Զ�~;��h]镫��%[�{�VnX����e5���EmQ#����$�:�]����<��OO'��3�������x��v��]��u��� Q��t��]*�Wo=��VE1]Mg�<ι�¦���e���9x� �������:W����-aփ� �ȧ���������+x��W���H�䒼2F��ۓ$1�m-_����r��}�4����{n#Z�4���"X��?��D�ced�On}����:z�'�F��>���ݶ�Me=�uD�v��u�ҽQL\����
�jZ�W�a���ߕ|�>ر����
Vfs��]���i��C��i���h��ԳD\�VZ�V�7k<?+4p��G*L�r,׺a��_�J�7%�L��نj�^��/ ��^#���W�9"Y�)cI9�z_v?B�w[M���x���}a��W��{�w����f�[���\�ekX���\�!�V�q�T e�(&����F_QijM�B���VU0���cP$<���<�0��$��c��(�v�ٳC�xZ),D ur�vSq#w?c3S_�{B��M�}a��k]��G=��;���{C��tOd����P'Nt�P���x��U��MkWH��6|�CP�m7N�Pd�.��߃-�S�:+���� ��W�J*�I섍����ċx�rƪ��d�)����O�����S/�釺��F�Kf�@e�C�*F��w��!�%�"X��9K�g���O�M'�� �߿7��v�Cܼ.��=;���&�����5���r��Դ�g.`8�
�9���ɢ�`�O�Ə�m3V��E��Y��-�J{	%h�#�޼�Ⱦ&H�R{$Up��W3}w�Q�W��գ�մ�wM�e��)Vxf�5?��x�DS(��p{�vV(��=�}���o��.��?���ݨjϨ�}1���u�Nc�#\�L2�I�#M>i����|�mA�"�<l�V�9E���;�zZ��=r�:�[��b���a �$��,�/���� v���mch�8��MV[���^�q��cv�[�5x����e�b�����7C�/p^㻁��ٿ�ޕ||~���#7�4�}#7;L��	�SCŔ�Xs`!|E��z^rf��4߃=��Fߦ��z�[����J�y���6�0��#G&I% 1~�Ь|_�uu]r����,�u4�R���L��ʌ�^�9h���y�yf�'�l�ߺN�av��O��t7�};��@ۯN��u���I����� M�pWy� ܣ�r�1m��ո5�_�M�)_C�Q���lW`D�����U���T�9a)=����u$��h�h�;mW��V�7�&�7_c���� p�x��k�om�ް��#��oe=�wc�Y��6����-#���*X�/���Jdc�6_������5�N(�q�B����hZ�J�cvf�f��O+<��H���JJ���a��%O�r��^��}�=>�-�z�3%�c+YC���_4�h�Y��*�Eh�
��}�����춣��E�w��Ӻ7p5,>��}��[t�b>��t&��9:vn|3��D}N��4�c��W�b��ށ�|m87&�N�Zƹ�|K,fȥU󽅒"�v�H��(��{,����� �~�kn_}FMA�BF
���	�a�7H����8!��8�:ɚ%�^����Mՙ��K�ݳ�2�:s����>�Դ�k����C�Ǩ�zo�r�i��q�LE���HiIB;�� ���Ι��ZU~ЩJ*VGw'�%@� �� ����||.t{jՋE���Oub&�Ӭܒ�B �$��*����������G:O��:��oJ�� E��}:�}=ڭ�t}?S�gR�e�ӾM#N�{���.���Ǯ%�)��U�+�u|��5]WV�q^�z�QMkW��N����AU����\�-�r��̋H��Q��m�3��-"��N�<�E�C ��IT( ���v�8���I�'�3����P����,;���:3�.GR�J�n��Vִ.��f�F�+�j/���eJ?��%BzSN�՚2�׋�ڤ$@��*<~>�}� $����3:�[
�ena�BXyp�S�Owi�����~�:�?H[�����{��L�R�y�zN����+����+��O�z{$�v���>"��hxi�<0�r��E<�?�;s �s��ۺF�Y���	Ϲ���ȣ ��f�4�wP
��{G��x�
=�^u���^���GT�z�P�.��}[\�����Z����;=��ܧg��v��N�8�*���VfrI���@ = >� � 2�*��E
���?~R$�'�ur�@?��?  �����ϯA�>�w9��%�<�h��6������ ��ٿ�����<��3�{��m���$�C!G$c��@;lPρ����� �x���� O�s������1"��T�͊_��UW����7� ��|�_�}��?��3�G�� \�H��k��A�;�Pw���������|������}������R�Mk��1�z�>�Ӵvd�N��\z�䞆ӯ��p� ���@S���(�q!-�_��u_]���h�[n"M�_�V-�׉��?5(�H�C2ȭ�#ǝL�^��QM5ccX�Qڬ�/�"����*,jZw�##��~�}�{1�_nGO�靚=��qtP��n���6��u�4�u�.���Դ�kk�D�*X�͓L��ee�����5z�>ږ6oO쩫<�#�U5�J��VUwﲪ�]D�̽� ރn].^�����PL������b�z|�"��J��jJ"�o٭4���{+�����u��/��}��1���Ft����6�Q���a���z2�jYL��l���Bn��޵� [�v˒�:q��e� �澚�)I�{�f�s����Q�bG�xF���K���yCر�2v�w5���$Q��M&B��3�,]���Gv�ɲ]��x�J蚝*&��q�*�4D2�������hd�Cn�B�n$���"K��FbIbI$��$�d��$��'7	@UUU� 
 
�z@� p�  Y�VB��k��sQ�r��_����6���̚��lO���� K-yx��j�T����tZ����b91��<�1��*S��<A�i�(Ixՙ8�e�m��^*����E%��X�"h�T�Qd�P��� ��0�,�DG*���/�˸.�������v*�La|��pm�%�i�=7Q�9���o�=�A;��Vc#����[pgb���ǉ0FG���"�Y�m��^�,��d���ߋT`	�����7�K�>}1�����f�0[kLQ���f+N%�b�B�}1�phEX���*Y�Q��6�P�,6 +%�;2�Di*����u�E<�D�Y��P��`F��X�̆����`l� B��2�g�:�5j�M�$�x����+QDKx^)v{V�����ZL#`�[�No�n�=�P����f��+`���0[ȪR�~���>m�<�r�8j^�V�4X�<���×!��C��!U��R8+q]�s�`(ȓVC�*y
�}�m�ر�W�UUc�� *U� lep����� ��}��������S�I����{?�B������8�Ld�qT�<�*�M1��B�)�Q�A;p,��S�K�ٹm5F�����2�� ;Y]@�0ۓ�b�Wf0�VSNs6e�,#!&	6�2YUY�wz�e!��}Xƺ��e���1ȇ��rV�w?�)��������A����9dE�Ҕ��+��V�K�����1��J���l�>	�S�4ځx���w�_�Yy�rQX��F6ޕ�5X������^5 ��l(sLc
Fk��*�ZH�:��xШ�`�����H��8dJ�[�=�D�U��L	QFD݊n���ጤ�N�R,x�7���."�zG�[}�Ȁ���N��G�Y,P�����c�M����c�<��;� kK֙w�tN�LSq� � K�[�z��\�-ma7�%�+�#<��\YB ̤��(�pX�Õd�f���d�|j]�;�� GP��n�=S�������Y�S� ����ȩ '�b�������[<�#4C7����}�ǀ9.��ے��1�V�(Q��'4�
��2j���8�À��0ӌ�2�0��J�QR��I�������(�;1��(+��g�ذp����䛒�a��A��"Q9�gwQTf�4]��
�р��*����ܐM/��i�n*�=Y��e�Uq�*>W�z�lW�q��K"8��7$�dTn�E�
J�+���d�&�y�7�PV*��'`x�VK<�X��X;�eU�jJR���5 �&�dF*P��������͓���K����m���a�T!Y_�57d �]�gw��"��JL��;l��4ē^���%ʐ��c����~J����U���(�?�x�O��W��L`r"��Rti��2�`B�-d��N��|��H��0�'r<�E5X��<B�4�z�\Y�x�/��Pܹ��Z����*�e�zMh�Ip5��B-�ёx�+��;��0(�y�!����c��o��Z�f�Im��G�q?f1�j��Ȗ=�_ʝIB����^J��A��,a_d��J(��
c�y�Ih�!�a�}�� �N�錷�(+YL�B���aIo�u��ߔ÷�'��!Ib�M��\b<0KcJ���
sf�3�2��Ǘ�bv�1����>�?�������N|t�	�U&�2^%}1�k?�_(8�H�Tu|��֯��R��6bY��x� ,IB�k�^��O��@0t���N5r2��cZ#e��9�)tp��E>Z|����ﯴ����Q���Ӎ(q��2���f@���(2*��g3���f�K�n��l�z^�;6>ƮJ�����*���R�7C-Q+�� q,y�c4ë4��Ӟ�yrd8TY�̌��:�]�nK�f@C�^,I�1�k�����Z��c��M�=3�#S�e��ڠ���<�w�N[���*�Ab�m�4���]ڱ�B����� ϧY���y�|��~D��?<�p]��ͻ�d��\���ŧ�MV�^���'l�>�Բ���XF=�����Kҽ� Ѵ̞���z3]���Z�'��̅c,`szw[���8��-Fp��6�̥_cv���lں��5�H'L��$����ö+�|x�N�����;�dЕ�Ǝ��h�����3ƈA^oSR�P��;��Z��K�A�:ץ�O���G���b_��u�(�`�Y-ƴ�:N��8h�Ɣ˵7�-Cy=n���ڞ�Z��`YP+� �}�F?Q�ݹnٗ�3���D�o�6/��t�Gz�����h� �o�B�$1W-ݚ��jZ�[t�Ik���꾫�4�p��O|]gY������������ �+}D�6�U4mKU�����O?����y?�{�q��}���0����4�Fa{SG���P�'�k���}��}{B�I�o�2�/��z>���Ɲ�v�r#��z?�:'X����4�,��;a��f~p�۝O�-���W^qu� sk�S�O`�ĸ�^�5���_Rk2\��ډ�R,��� �Z���=��6����T�Z���Q�OeV��Z|��U����-�O�n��P�g{��K{���=��k^�k���׷�M{B���z��{Ӛ�V����u�v5n�״�w�y:��<��!��TL����,��q�-wU��O��AHۚ�p�WV�Ejz�-�4�%X���j�,{-SD��>�^h��z�X�X��DV!,b4����O4}��^^�I�Z�}�j^��.V�ܜ�/R��]��Kh��I�=W�?�b�WD���]p��>Oʎ!9WZ�*��I{H�.ݷ�TВ
�_-t�QY�q�� }~@D���<�5sY�onT�x�#O��3��C0V)�X�����` / ���_Q���/��[�WGc���{��}�]D-W���ؙ������|i]^���2kT�xf������+����v���Q�r�ʀ�`�s��
MT�^���`P��{@�q�/khW�k�OSe�t=VL�P����9�2,�?%�ƍ����>���toR�W�][T�u�<�G�4-G+J�1/�f��Դ��طC��7�����jT^���٫f0��*,�:��J� *����8 �'�}��vH��;xf��$WWeI#d!���B'�m6���v��>�����_�D��~�����,�NKM'+1 t�Z����y>�Q�M���
ԗ􍩤WԪ��|�J�h2�H�TY�{Io����]`�j�KV���;E#g�6�*v9 ���CD��r��(��� ����ܧa���j?�� Et� Uh��IW� Z���9�wO�o���6�ӱcj�m~�A�.Q�8�fQ�#�¿�-��j]K�)m��a�b�Y'��ba�Q-b� j��&1I���/�߅���=>�a�5��S�K��ib�fq�{?@�a8��F~�HoG|=�����������^�T�Oo:�q���~$�t��ǩzsK������<�6���m�=>N$Ϟ|3Żw�����Š5�5KF=J����Ӈ���W�?/$~�2��Ֆ7�FX���G��[WB�W6����F��S�&��0��%)�wH�B	�C�$i�&��������>��.�{N�+c���ס�k�3}�w2ȅo�}%�;e�_"x�֜���e�ѕb7�W�c�.�ٷ5�3�m\4��j��T�'֝u���',9��@"0&L��wp�wI��l�h+x�&�Ns���!^u=;���� �� ���!
�ӫ�c�^��7K��i;����>����Z�W����tf����>��8��||�&�:�z���3�t�غ���Ͽ�����N��SI�h���
W�J\��Z����9��%��IXv!ޏ����J�^����X�N)�[�,��ڛ�{�4�5c��C,S�@,|���ѿ�V�ٮ�����:�U�p�v��u��t�_wY�ɶ���j]=�˦t\6:sK7/R�`�+��s�t���Q����<Ӓ	+�q!K(A�p�q(��㙙�^S���d.��fT��c��6�a+��]�`����=��	n��}G�}�wCQ�^�{���ם����Ƿ?�� ԝXp�4l�GW�Ɇ�ލR�~Nr&l,*i&�/BWW�v�M��������Ƌ���N��H�\,����qخ̅;B<hI�]�w潳����|l�B���\���|��<���~0{e�e�2}���{K�~�{4�;�㢻���u���W�=˦��􎫢cj�Z����r�Z�i� 8@ǿ�X�:�<�P��f�֥���^>'����J�|�[� ���(k
�?���M4�^�;K^�$���wQގ��9|;��W,í�nM�%ֺ|���Yj�)ڲ���爖�k#��$x�U�n�� �Zw�ݗ�^��Gn5��@�?C��{���^ʞiYg��� ���ʦ3a�S�)����T��t��߱���䍣�'�%���g�H��8��H�#2�B��#b�����X�j��X���7�T�� Ep�Cid�ܲ7h��
��#ֳ�ۨ}�jx���^��ޝ�`:�W�Y���'�i�9�/Hfk���׵�:�G�.��q�(��CF�9�q1{)q���t7oh�r�����V���V:���]�Ŏ4o�x���SI�0�+#p�<��Z^7���ƃ�T�����G�/�=2�HuIyk<q��x"��a7j�ѯt^���b�z�g�ܮ��� z�t7�����^���ƛ��f!���zd�ok��X���zw�L��Z�|a����U�oi[�R��m��!�8i.�Y;��(X�|P��!�hsc�Jt�˸u��Jd��L4d؆��HU+4��KL�%������qע=����T����OpX>�pz碩�%�-o�5>��h=S��]g�m�>�����s22 ��L?Q��SL����UmBb.|�#�d� 
�K�Gk�_d�Vo]��7^I+Ȱ�\((��(r�r�U��K�>�,�<Ӹ��}��!�ۢ��1퍢�>�����Z}ۚ	j��<�|�غ�?O΋�ڎ�b>#������ݱ4'��;e,s��Ry0��L�~��/jI<��G=������ꉐ�$O�;9����.���J�d�C��^��s��0z_Q����+Q��qz����(�={�'�B:p\}N���`�m�~��Ab	��0푘�#���P� ��1�9�����RX ��0�{��{��%�׼�8�w�eZ�|��C��0o)~)�*F�K�1u]�r$��mй��^�$i#���h9!��� ����~�j�j���.���O}���$�\{�4׭N>���Z��6mV�Qǎ���;(Q��lϫ�V���N��� ��r�iYg�?�y� @��x�P��fVܙS�;;l�`�u� ;��?���(��e/۴���!H�$���o���>�����4��I�Uܳ/�+7f]�@?������ȱ����� ���R�� v?�?�)Αk�vc��r�Ħ>�ѝ¾	���`��0��4��U�Jr�/�9Bw�5s�&�\��&��A3	q���_��x��!����	�{�>������zKI�i���s��a`?6<' a*�G���+_���+��d�+��,�_�����]�ʁI������Y�SC����kؙmSO�O$t�����z��Y�PԤN~Ǐ��}����eϾ ��2�x�|� �y�~2n��0&��N���1�]��(
���Ăv?��bсbЫ���y�'���e��f��^~ ����={�� ��R88}C���!��I������S�Dm�(� �Un(,�u��W�$��T��z������e4F�)�NZʜ�H��9�_o�����j�Y��I[h6N��G�q�Z�@ǆ>k3p�>C������]΁�o��ºI	R�>�� �A�f^���{�\EZ'�{� ��g�8������s=��w�{��o_�o��Nt��ӭ�H�?q��ld��m�e!\��W�0eL��r�2Q��G�[iۋ_�I�]��w8��~F�5�w�T�#�U�n�Q~��Bʊú=�[�G�$mͭb;���D;�fِ�*Ӊ��{X���#?�J���'�ܯr�������s՞�;��7��^���tGAuj��L�b���l��Ύ^��c`$1��=+f�lT}[C�1,fm�׮�m����+�~�z��
[B�~n�fR�[���i�A-�Q�Fc�� #;�5�\�rG�v���#V�Vzֵ�ѷ<%�o6�rIxDz�J�����?������C���f��s�{�=k��K|}c�^�=�h:���k�i�>��\��kS���Fӳ�=G���d��:N#Ny����������g�z�G�n�~Ν<�G^��lIhF���b�`#�]mi�BEb(ţ��cu�ah�CK�vY:D�"��}J�ylQ��q|�G^�i�w!ϧ�5-@�H�E���v���h%�`tg�4��wG�aݭT��n��s����E����/�>�ꓮ�ܞ����퉁���:^�?P��+�m=$N�l~������xi�hۇii��i��n�"���k:�Đ�J�d�O4r<vlJ�⊼\���M鴺����<�H�sՅ,�W�k-��ŧ�"F�ٔ�a#5ብ�I�Q�����������J�H���>��~鮒�t��r�ӧT���oLh<������sa�>�0�6�Obg�����|����}��=t���w���[S��R���U���_L���}:��=��T���2 ���n.�u#V�j�z�ghi�ㆋط37HlE���=�r��G��Əus;���Y�g��:Wz}��k�η��ھ��GJ��}{���Y��������c�+U� k���:x�L�z�|�7�_	���.�'Z>w�SK�5���{-���T	d�& JK,6iH�'�X�J�z;�/@����VԖFӑcI`orV�I$�BY�W��d�,Cf5Aђ��O{��{4�� ��k~�:˾��}�{Ҟ�ڻu?Uv�sКF��OU��9����P�� �E��Z���r���V-��_�����﫚���6��j��iU�:{#��������k㊹r�us��G����z��sUY�UIT�Y//���N����߻�!X�r�J���n�3�����폱���,,mW��� Qcj:�>6UD��W\�f�]�^\y[��!{����� Ǟ��5g����b��e��W�b�'��U�VP�������ȧЌ4o��ǭh;o^��G���\�kBB�P�i��2���E_�R��=/鮌��l]���:���o]���>��gq;-�OX�c�k:^�������<GDˋ��W�1�F����hC��<���6��n]#Y;3_����V܍=�`����$a�@)k���9��z{����ݬ�-�m�t>ْ�ʨ���>��ڭ?��O*I �+��Kg��b�ĺ��]C��M�W^�빝;�hٝi�n������vl����tV�������`�x$�B�dM��L�u=�<����X�Y ��O-s��qG��g���Bs,c��[~�Yû"mLJ�{��)�+���+ۖIfp����1�Ԗ ���^�~���{-���{�^�w������:(�~���k������:n���V��V���ة)��-h�m�ܿ�~ʷGAӴ�R�:�r{Y�$�+��0�����/�V��;�=K^�wT�u�{MLT��SN�4��n�q���` A�wl�\� �/m5>��篻k�K���?g�{����}.8y�t+g�b�둊j؏��lI��6�'
��w�1�����O�V��������9F���)�7i��;2�
�%]d�y�9X��x��ܿ���ǡj��if�หR� ?���{$=�#�QD�2 c#v��w�퇸=kߏm��1�m�m7�0���u�\u7\ai���c��WFjAl�_QZN (�8��x��ǛW�?��ON��>�u��{%5�s�9M��hӕH,H�,Ĝ�_���w6����M����
��ܨ�Щ��K3w9��}l}!�_��k��GH{��G{����~�z����;K��m95��k�xZ�5KU\*����u-�L5F��ʩ6�G��m/��"�]:��0ҫ�-i�Z�5v���Dq����'qv=�F
�Y��e�������5MW[�u[`Z��*qXE��o"��Y<�:�
P�y":��f��׺����x��K�z#/���ֺ��)��kq��8h�zn.z�S ��5����D�4b�;��{.���tM>�2-Cz:sCb1v�D3:�!�M/gk!�+���6wDvN�t��j�W��z�ZJOue�D�s�4���č!Uu��g��܇GkC���gvi��:�L�9a5�K��mGMְ��_B�W�ItߞN����{��C��d��#�u�/I�Ue�"�2�� �:+�e"��r�Ϯ�2��:��$3�<���U-��S�1����x����g�;����zש��h���헷}=׽e��E������Gbu6���wH难KC����W"zgK~&FE�SR��w�)��t��O`F�P�(�s�m9@�݁��pr�i��j5���y-(����2F䏸~��f��� ����=�Tv�o�twhu%]'�:�'�����^���۪4�����-���7#�t��u�iMS+.q��Ʊ���a]UX�^�yd�1,�O����P*=��H�'b�H 	$J@����	���EY��$ v�G�_�����v�ˏ���~�rߩ� ��X��nvH]�o��� ?�����G~?��� ,�o`� ���v ���K1j ����|��ס����椃��i̓�]�n	#� �e;��� ������?o�� �?\���=�����2�8�3Q��a�7�� �#�� >�#�������L�����,#$BնS��!%]�j�uT���̪���g1�	$���$�@ �< ?9���ʈ�p �I� >�� w9�od^�1���=g����`매�jt�OEi}5m����D��>�K�m�AW����d��T��c���]�ٝ���к���T��ؖi�mN�)r�dx�
�^.9W����'9��v�֨ږ�x��9>V^��U�Dh"~�V)����ʡ[ꣳ���7�>�ew{�]�]W�4>��t���tu��ei}7���G�.�O^�{hJK-?Mӥ+d�*��R�qu2���_J��A���Zt�i�!�V��U"�f'�ܽ��HU��k,�.�&��Ff�wn��I33IfI8�AL9ixT��2��2�*8����p�n�е>���u�'����u�mx�=S3u||����:PR���|y�Qh)_��77U�-B	t��L�0+%�Bԋ�R���V_L���$T><���h�u�u�Ω��U��^Y�B��۶������B@ha2~�9��~��=��D��Q�����ǾNC�^Ik9��t��+,Z*�g��qZp�"<���I<���9����7HÅb���ͱ�[8�����2T��pȺ8�o���R��H�8��d�G��3� �y���YF�y�8���ԄԴ�r��"c�_"�o ��@b�,>�����64��M&��*-�s�98��$�-�T0���s�8�!ڮs��@��j|�`�Hp��`H���zP�jJ�6`�y�>�<�@��?�(S�ʱ�G0L���l�� 21�1H��������Ϳ�H٘���f�E&�#�
�w-�(�7%���#|LayP!QI�d�5�M����+�.���(�4I�7���R��i��%�se-�������m�ܟLb�շ�p�f����H:��:�����;�����c>J�Y����u2y��1�HpUm����T���O1���90���� t�PQN���ǳp��*��yD��53��Ce-2M]J�EY�� �����1�2n*l�j�	7�p
�v���lF��k+����h+|F��b���q_����v�X�X�@'zx�[��]��UI�C�L��r�0�G���6��\�X�M�'v!?����s����yA7n@JG�y��eM�w
ۋU@3UR�/˚7�Ldk� ]M�G�)�3����+H�!~�dq�g�a�R,ʏ,�صy�(�9;�q�8�	�,�^,JHe�2��f�W��o_�����qqm� 6'����X�f��q�'Ί(�X��H�(g�d�nY��B O�0N�Ѭ,�gǳl�8�u|N������w*����(� ^W@���q��Kq.�l�X2��@�8��H-錡�vo!��I��]�B���Bȹ o� ����1VP���V��IɥT������I�E���'��5���TUkNʳy�	�*>:�m�u���uc+��U�/3s!d�MԄ� �^<��q���2_�.�Xҩ���1D�����b�_�)�S=��vdd��M����k�N,��B�R'����#���>r��_"d)����w4�)
��w<�uc�w�^OX�K��[�SrU���
�`�wPx���z����fne�vY<V��~]�	gn%�,d���Ab�K~�� ٙ����X v*�X�/(��T���R�)Vm�3fH*�T&�zU�ޘʛ�%���چ���i�lV�N��\�� �#���0iO���}�QK�(ZSU!q��ep�-ǉ�zU��7(�+&?+d$Q�ݖ5N!8�M��nc#-����`����R��RϒUxoȕU⨥��c'K��Th��vE!�Y'96��~L���y@PH�� �|��fe1\��F4񙯑ܝ�&��.�"�Cj ����Z�H?�@��#M�~A,b�R�����-���:ѹ S1͹}��F�zc h�J*��pD�q>;Ys�21g��d�U�7c<�k��Ɛ�%�Ɖ'�*@_����Ɋ�i0P��Ix� /y��1ٓd6w���H�c���h���Q�ǉ2�f-1w�R�C��!�Ö��
,f����J���9(O�RU�=B��>�,X"LR��'[Џ���� ���m�
���=���Ĥ���V��Y��4��vc?�rI�T�~'��h��+5Ւ�
��)1����U	=�)� �~E��I̞+vef	�bU'Lv<Ԋ����RĮ��$ >���Ґ���HL�e�CGV�]�i���� 'pU@>� Dbe�֭*��RkW�g��lh�h?o� 31�3%�ERoe�T9j��9�QG>ly����6�d�$��lr�rΕ�p��o�t*Qғb���+��U�c<T�v6�3�X����b��2`��jf�t�g���h6RX�9��]7[���|ީk��B�J%�q&�|qE�N�V�AZ�MwU
�rW��ӝc�$1_#8~nU^8^���Er��iX�^�E�!_���r�;=��Z�7�]=�k�T��嚢���9��O!�O�<���B�LgD=�wL�mQq�MSM����rc4���/-��h8sU���	@��� �T�<G؂=�?{�� A�� � ��z �#���+��Ii���zsKP��ҳ21s�t�Osl���u�-<��>d�&c]��c�i����i�;�˸��Od� K����G� �x���|�s�7
tϭ�c|A�k�9h6>𲒙`
��m/%���jN[�KUTF�5w�6w��G�~�aiy?�:&�L�2cag�'�䶢���3�ѵa���ɍe��+� �-ޥ���$n-��Ŭ�r�hX:���"7�>J�ƾ��H��2�K�m���ߺ<�Cw"�D3D�I�l�2��.	=y_�ۑ��>�{�퇺�[�Wn������];�w��pt�CN�]h��1�c�g�����uM;7#?G&z�?!pz
a+tg�6��{��EV�fM6I�Fj6�yf�i�",QWi�8�K܏ZF���e�}B��n�U�vک���zUaԍj��v�ub�Q�F$y,�����l�b(��J���v���W��^���z��g�
i�:N��X� N������M���ڗMu�. E�6V\p�D�g&iMI����K��=�5-C�,����JһSH-V����ɧؚulȡL�R�r�3}y���ˣ��A��o�v��=;~[Q[*��sJڝ4hf�$%�;q�I�,��hBo����U����o���������OI��Z��DW)���135�hC�n��.~��E��i����Z�w��}.���H#�{�,ī�n��A�3����)�n�H�D���܏|�Z�G#�ۀ����m7���{�u�'�� c�^�vwDN���Ji��6GKL4�����*=t���6NV[~^Iɥj��;��/���:���w�C=�,��t���)��rٝ��&��(��8�? ,��|�N�v�N��~�I ���_�	d�FK��	��(FH�T�O1� ��>��O�����t��ܮ��OC��Om;W��Jc�6�Ϛr�(�j �:����1d,1����2���|ko��:BM��N�\���̖fh+�ЎE���:�)���9�;�6f��ZĻ�JϬi�W�E��^9f)j������ ��B�C��x�����,>��� �~��v��O��{�����?/�:]�5�q5s`�阱E�=#�N��c���k�m۹��э3bv�ĵe��R�ē��"�!Va*F��C�><����n��6�1�w� �޿���Z�`N!
���^I@��ܪ���=P�u7�/w}a��z�Y�Hb����n��kO�:�V���t�{N�ԟ�8�_�#
��<����~��wR�cKW�E�m�'�)��4u�nȥ�W@���yvB��;P��+|D�-k��N���I�CY��j�:sH�{3e�x�n�(x^�����/a�ʗ�O|���}�뚷P�]{T龛�.v��h�]e0�t���n�z>F���s����Ȅҁ������[e�p��}Hi�A
X���O�P-:���5<3��#��/r,�������[��N���h/���b&�?0��*�o��� ������/�~�u����c��O�����}9ҽ��M[���X��7M�]e�z��cCp�Y�X�����ό�p}�����:��>ڒ�IbAV��	��)�c.�"Q+����V�J2��{[�����u����Y���mC7�Q)� 1��q�dXHA���ϻ�N�wg�;[�]�w�;��SE���`�kS7�t��b� T�:{YҰ�S�^��-n�9u"*��hy��tK�m������-Q�riSq�k��
a��VwHnR�`<�:2�Z85�G7���+[Cr�z>��_y�:�r�H��^H����n4�G�ܱ)!*ܪI:�s��z����]����^�h}!�jz\;�틻�Z���M��Y�n���OPՃ�wk�!NuS�S��3.reɷf���vn��4}nX"��;�IX���io׋�]:�s���
��{����7R�r��iͭm0g�j{sW{
�:�i֤-� �#y8�v:9X�_���� �_S����n���� n�ރњOEˢ���:*ݻ�	cW�/���y�k�����~9YCRŞ���?��m�yW�GY�n�J�*���a��	)��(X��ȞTs+L%I�%y!uh�p|}1طz?&֠��u��+\[1Xs0f�F"h�*,F2|,�K��w�ޮ��ǵ=Yڭ�:���nz+Lӻ��X��7^��Pt�\�?K���ֺ��eJ�41��f�q7�m��͵�i}`�dҵ��	� Z��
�h�^�j����`c%(�]W�--��׹{�WO�4�rI@NT���r�ȐJ�򰍣IO����I�,�lK���?�w�3�:�V��9v�5?n]֮.T22?^����]O:d��i`:��ц���������t��W��B �I�\��Ԁ yBU�#�i9�Q���<�[�N�{_���y�Q��E��M�c ��V^֞�xK �摤�C�{�#�>�{Y�;��}��;Wڞ�{u�������hz����9�Y�v��� �3�Uɠ4�XU�Dh���./�P���;c}7PtM�Fg��~�4b��k=i�ĝ�d�FVY�+3�=r�{dV�o���J���6��E(nmmU�D#�Vj���ʃ�+#���/*v���7����G��ֶW{�:�ydhQ��w\h�v_�m.���^V��<����v��l��U���8�u0Zb;~b>�~<�r�i�b���l���f�ޣy4Ⰳ��ܬ_��G-]���G�3���_M~�=����p]����w_�4<n��^��������t�5�WwO@�Ý���$��2�.�B�@\���x�z�4��+&��0����{����4�� ������+e�>r0Ƈ�L��Ge�,@ p��nI�W��{�'5������_T��׫:��F~zit����HƵ8h�^�)i�V���v,㉊��8�ݚ�rM9��%���/ط'��rIX�O���E�梹$n�j�n9��d1���_q�<G+K�z�r�l6��.�͉�)��	
V�YoWP����ubwPw�;�ڴPW�pX�kKT#F��yVN�G��pO�3 ӥ�H!j�yRs"�ʆQ�����y� ���u&��3'���O����ӕ�����r(�R0f��n��]ʶ�g��W���w،��!��2��%��a�X��mҊ��3 �?�x+����+���4��Z��i�hY�2��eae��~��R����8�x����Z�:21�v���G'�������e�b~++�����G�?�?L�Z��Eֈ�L��)��� ��?�� ����*L�S���^����Y��ڞ�j�lv8�˨�bc"�^��2@��� ? ��Tir���G�S�x̏���Z�>��
屔�V� ^t��3�-#�ᆳf�5-���W�n�aD�B��$}p9 y�~��_����x�ȃ�����>�� 3��~���д�f:�Nuց������Zݫ�èi������+���f�S��%�^z��ߎq�Z^lޚ�j�V����g_���n���A�6$��|n���Ϫ/���'�2��y ^��"��O ��x��J��u�M̄m�����Ĝ�0Ni�1�e���ъ��� -3���ێW�v0��
~�?O����·2Q��}}��!�0��������79x���o��/@m�XzyK� 0m���XlF���.x|������ ,��Y�v�)A�!O���� /��M�u$�aln���|�9GP̻i�`���Q�L�
I?*w�o��'pi֔��>K��>�Oc� />���?�3 Ү@{�����9+�������{ޜ��w,-s���멵����g��sU�:�\��s.�dt�&|����cO���t� X�]��5M^���Y�+�]��F���G����ơ�G$*�$�����Q�n槪�,P���珲���B��}��Χv�GazW�����vG����L���n�ԝ��%����������o���]QӰ	�s�u�u�Q��$t��:�H8͓�m�-�CD���j�O�&y����fJ�(�a,�~j��H�MY�W�!�K0:�H kڞ�f�M#m��c��'�
Moά����8�M>�NS�+ʦT�b�N���^�t�f���~�tn~��/n�U���C�������;��m�,O+���֥L�#��9da�uWNWX�j[���'��67X:G��}�f�Zƙ�Gvӯ�oo�x�hV
7���Zg[1���W�!f��^��ޖ^��f��X�t��ԧ��K���Wф�B�e� �oO�#�y5-4��+�8׽W�vo�w����e��q}��S��vwD�0�z��O�^��^��~���fd����ۜ.�͞���	��|i0��Գ�:&�h��	G��t�M�
�F7k�V9M�r�N4�yݦ�8�~�]�q�|wȫʍ�պ�����L��U��7�d���߻H^d�w��F�9�-�;��q�g�~�;�;S�}��p�OI~��кKP���r�,Hi���A�׳:?����ON�������̸�m��[N�|7�Cܚ&���l-ۺ)�Z��GVݍ-�/׍l�*�xS;��N	>RI� �,e#�ځ{nܻ����д�-G�<J�/|0S��Q5�hY"�M;��V"�uAV$%��gW��%��wh}���ٺ���fv�J��i���~�v稴jtv�L��_+�k�c�tA�X_Wh�=s>��Oi��?Iw7FzI�!Mݫ�5��l�Q�Rt�ߨ0E5�l+!�9�+ ��`�����ZQ�����G[����R���X)Y*�w)��cYY|O?2w�C�g��{�ߝcܯI~����zW�����C�5.�h]m�߾�Ӻ�<j��������԰M�1�3n��\LINm<^5���U��3ӱ����U��&V$;~�Ib���(��0	d�7jo}�·.ޤ�p���U�<d@�c����%c�ξ+,Y�d��'4{����j}���A��O�{c�^�i=��{��w�K�Z�e��g.��j��y�W��c�T�l�l�ŒP�Ύ6��Ӊ�uO[iw6�����ф�f�P�K�cb_"��k#�������?{�X��D��v�&������I,�=�(G�Q�*�^��H�+�2�A�;{�����{��L��wU�?�Z7Wj��~�Mw
��%m_R�m*0sg�%��K����}_⇥�M�����j�:m�Vz�4�B�� �B��<�����%(����9GW�ǩ{Vз&��i�ͽ��X|�.�'��xTʮ;��c++s8;���ײ����}�'~����>�=�ŧo%՚}��аtm2=)�:�d0�d�f��N�0�K�p�,�n]﯄]�.ﵨ��{�n dj�C� Q�
-��B�*���"r�)��#��G�6�}R��p�m�&i��hwi�rJ#�)�]ۇ��)N�H3�w{=՞�c�ߴ�m/�+�^���w_�Z���k�\���~��.�u�TNP�r��8a���E��>m�7w�5�Q���Q��xKK���V17#�;��Q�F��s\:���_5�Z�CF�g�����h�J�(Ҭq3�х����u�#�{1�� ��^��^����?p��а��r{{�}q�k�OV�mCN�L-�'�8�4v�$���/<�m�d�E��'z֫�xc�uh�L�UX�Gv��q�F����S�Z������e#��{z|��4�0x��Yx��uڤ�v�����[�������}S��i������N����ZvG��}&=X�+�j��315KW�Mz��Lq������D���u�/L�;�����#Ա�j?4��F�Cj��3�;�,�h&(YeBT���7��}��ۻ�D���&Ts��*�X$��!YFLR4�1(�H=���WF�w��ݝ�:�������p�Q���=S�t~���_�:�_�������D�F�����Ĉi��]�z��s�u����r	��h�r��A�X�x�r��V8�(�݋v�cN�|3�6z�]���غ0�
��"W��dD���Yde^~�q�i�|�
��랊�?P��O�����0:G�u�:K��2�>��.���V�1�S�[V��*6FG�>J�J���w\����t�LU�c��Z���iA2FaY�� �X�S����G���N��t���=kW���y+�8����%je|�G�iGwC�3M}�{��y����_bz�zc�Gczy���8=����e��:T�쌽b���}3�zs�2�4��|���o޺���[� S���H�u�bİ��l
fvV��+ �,�I��7�W����Gg�/fɹg֍8"�I�m`+��[��
Ȼ��d ��w|��>�;[��� �{E��u6gq�.�hZ캻;�q���uQ�Eմss�����M�o���G�L�`j/1j�*�5&+�k <,
�Yʕ)�!J�a˃�2����,�����%e�`<%8!�>�{^Ga��nD���o��K�kZ����c�wf�WV�Ϸ}5��9X�3�B�� c��<2/)n�t�L�c׾B�cG�8u�U����0���@I�E��/yv����)#<��C��KǱ,O�;��w}����}�=��i1��'�\N��oGc[G��Ea�#+"�Ӵu}�.����ʶ~���;6�4giE�t`G-RV�=�5<���w<�� /�Tg��1�9�]�	�G���}<���,}��U�QbJ�;��I����o� ������O�}��� ,(Th���R�)��EsW���t!v����};y���p��� ��~~x#-��@m�!���9��/�M���m� ��� x�s쟱��� _���KЀۧ!��)Q�܆�r�s�?�����_��>}�y� \~?���]�TSmߊ����wؒ;�>7�_�����?�~��~?�.Z~�}W�Y��.N�Ǖi���m@�a��ǟ7!9�&�WMC�w�KE�(����vCc�s��O'�UU�؅E������T���v��V� v>�>���.�Ҫ��}('�;�����5_��Gw�Z���֣�����t�Yv�X��?����hu��]C���o��^�pst��c�N]���v�H)ꧨ;{O�{�^	4�>c����w}��#)4�	���5�hY��Z���zvؚ���a2�f�+̧����́�oq��@��q)P�֏p]����o���c�zdr��2z'�9���^�j>Q��m����|���'U�+Imf�yY�1�Cz_� �s�}RS�]���@g8j�m_Q$q�F+�^/FiK�-�gn�SR��m:+Wk�<��|5��1O�Π9$b�U��"H���H�s>���5�͞��:�ڮ��N7At6 %&�� ����o�Բ�dY�BK��#��K:��,���#n���_�ǡ5�Hb~>��G��k�2���kh���Lu=fD�{N�
�<�*�%Z�� �FK�@{J��ð~�u��Րe`S'�zb$1�c+�0�]U�,����EQ�$4�l��̛>����v�������D8S}2Ch��V��Ȗ�HM|�iF,���B�n����O�1��ў��-�וb��[,���dV}�C�K����hX5x��>2!�̍2������V1��I������(ҩZ#�t�����j�GŘ��c�
��� ��O�IŪ��ugW����ɍF�6D�6�1�q�q>�V�G�w�v[I�t x~���پ 9c����c��	i���T/"���y��3���C�܂X���$��A.�q�N;�4�ȧ���$)��&��LdТ�U{���HK�\���G���E ɋx�&��@~�I8q|�G�t�`����z�<�r
_�OϦ1��@�u[Z��
�8ř������`Y�b9|��)����8�d�fJQ߃Ro!�;L�^Le9�6@�/.v��e��ud6���s�p$���ޘ�n8	o��M£�Jۚ���Sa�; RT�� ��2:�%���l�eG�AD=1�����*Sf �G�1��Qx��4�i��<O���3ȫ���v�o�ԍ_v�cp�$� f|E[�RZꦇ�7�O��.3B���⁜�M��@XI�� ��;.��лrc"�+n��� �',m� ��'o��� ���Iy�y�ў�IcxӅV`����E~\y8��R��2�!�*�+�v�	0%\1;Jp�c"� l��F���c���L�;&S<N�,��Ï�t�
�)UL���<t*_�P O�l��y7�1h$��e�r�
yL��o��(���r9�q��v��U�Hxٕ������Mj?lT��f��ط.J�Ic���Ug���h��u�[p�
�mو, !QC�TVN��6nfU���ɻ�RS���͸'O��c{���Ͷ���M5W�{.��%�����2�R�TW_r̐3L�J��IP�L�%w�AV�6c�2�{-s����eFSg*���8r<x�E,97�1��g$��{���Q}����r�Wwv��̾G64��Fd>ȴQ�Ҙ����bJE�J� ��$�P��'>8��Us�!��T�2Tb���>���ֳ2[(	T��o"|
��˪��8	�V;��%�Q�<V�Wˏ�;���ƒ��S�$
��1���3i�lԢ�U%+HI�U�$���(��� �����tje�6H78ԩZ�rEE�^d�m��\+r� o�1�Ǣu*��
�[��uP��I���rY��Y��X(c(:�Ʊ�M����s�:�����rpW��2LdT'���N�+F�Y�m��a>K�A݋|�0a_�z�eFb�'&�9���9<R��((���3�cf�JГ�s��il���dUTa�[nS��R�Lsjҕ��"�p�f�
�=�Ven~J' }1����UR�u�jӫ���Ǒ]�ɑ��y��G�~�aZ����Wʣ$��J�]�-��l�g�4�!�wb�@YY(�R�(da���0��]���8�c:E9"�L橊�Bd:�5Rl�.���[i��n\�Y����¼�8�
����Q�x���%��*���K�(]�s�2�Œ!k9�&rU���f�O��ķ9컦���1�i%��/�M 4@˿�u��yԭQ�'� �0h�`8�W��v2At��t�^~
?8�E��fIL�/	rM҄�v��b%2g�c$L�-x'#�����ي�;�>��%q��H�xiN���G�L�����I���b�	y<�g�*��V�I���Ho'8�rY B�C�'In�rx�� �آ���W��Vse,'���1��Sb��ieb�)?�d��WV�dJ�dT�n_�b��@b�d:Ef2`Ւ-�H��Z.C����+T�X#���2c��x��g�����v���L֧)�VT��*��1��fy�zщ�[x�$��<$RA��E�}Y~�,g�Դ_�
22V|'Hll5�5n�=���Ϳ�3yh4oLf �N���-��RVJ�.,il��sY�m� 1wA�%@vB7�3C���Mֳ3뇦�Ʈe��������?b�/A��1�(f�Y%[�����s'�^ڵ^�}C3�c���o��@�X6N>.4���h��ğ�J�����O_BL�9Zz�5q�-s�NFE��4`�L� b�:��g��}�}��ez�=[�>����O&4�.A��3��� �GL�����^j]B�u��m-�v>�ږ��Z����a�j?�V���2���x��a���C��?�=�ǫS���9�,Ԙ{[��U��W��b �]yS���y��]��vOj���hݲ�R_@�^���[��|<x��o~>�3�^�e�'��#�2���A����v��G�Z�+��=��%�'<��a��{LRJ�FDZv��](��=��f�����5�t���vޯ\qn �[�jB;X���:�ޏo]�LS�X����1i�F��3+X��]KO�	uy+42��XeV{'���?X���)��𾩤BB�e��?c��뀼>݃����=C�&��6k���]����A�� 
$ ��Hc븞�`u�e:��5�M#_����jX�P��U��Z�����"d�>6BʼWps�&���6�oi�ê0�P{I
A�x��^G>���׶���5���j<7i��������ݿK>����������L��m:cE����� ����z�\��p�噤�N�-)1�4���S翑��'5����.2Z� ���n� ��)���u,jd؆�d�)�]��8����8��ǐ��{�:�F�	�<���UЩR�4��R]zp���|�%����)D��v��4'��և�C�-R��T���n��.����wM��wEi�]���ǧͱ��s�z_*W�!��r㍓�tf+d��:��z��&�Ե7���i���z��%�ҙ&��H����Ī�$�#deh��G�{G���ޡRӪɹ�mXu.Q'Kkk0�R��X�Va��B��I8])�� Y��c�v_Oשz��:�V��3����̪x|:~��q�2h��~E��M�	�b}M-|�:^�ZE=���kq�g�f�*�_@���G#��נ҄QדT��F��U��Tf<���䴪~�e1 ��;�N��=�{�>�v#�;�ޮ��?Pw��� Eө4��f��Y9�r���z�д�}K骘�S\�z�֏iL�s�3�����N�-�h�d��B������^��d��q[���ȑ��EpU�G�}�vWRt*���mopӎ���J�]�bG�NT�֣&�%g$
]Ǹ�}}�{H�Gq}��r����}��/Pv������4����iƑ��A�����e���'TFXF���}e����٧N�)Ρ^���i奨G7gsE��ȏ�J�����_ze����i���*�R�4�L?1��~����V#��S���#��_��w�F�l�������~��4�^��R���+�zfi:N^���i�jR��yy+f��Yt��m+ڬ:����s��85�CS��K<R/q��ZTT8ۂs��\�����ۛ���H�~r��=���d�����H��OҾ�u'؇Pu}�������u�={�g�A]T����>.~�*��n�����+���?>>&��)O$�3h?�v��M�b:kO�Xѫ�^J0$~X�I�e�,u�X�m耊�%�����}���������E�js�b-Nn��i��0�D�;H�CnC���d.�FAe���~Q��u7u�P>�f���_J�f���w#����[�׺v��cc7H��KK�]9�[Yʍ�O�x�1u���SP�O����e�b������O���<����;H}�O=�$ỎnWS�]��T�ۮ��+4Q�[U�eV&i�t�"�O�f�d�T�WTq�����\�{m�/�����S\�%��s���~����hx:�V��y����+񻳠�#de�O7Ư�T�y�P�غnץ�����z��C_������Ka�Y,�9d~�6p�����.��5��{�qj�����+[ն��2i����(+$�k4�P���{]�����V ���w�=�t�n{��y���.��[t��W����.�����qմ
����o���/Sn"���@eΚ����mן�� �w��hޥrA#Ih4/$6�t��-yUB$�&��
�l�F�����ߺ�n��S0Km^d����Vj�Z�X4l�[�@q������{{����݄5�u]�|�m9��R��zK��]^�&|pzk��.�?4ꫨ6�듋,<2e�7��v�Κ�꽝T�ܚ]���iR���}��+�i���፞��~�Gs��t��"�e붫�ƜV!to ,l����ą�����߫^���{;�ߢ���i}������w]�S���:�ۆ���`gjq���/���y�fŴ�H�B��.��7z_��{R��j�����ʑ�YRc�[cuDU'��t�]��!%FDfi�t�=7��_W�t
��ޚn+}�*8�}1�FO5����v��{đQĎ(�2��{i�lKI.ؼ�YMҎ9�A�K��R>�������ǣ�>��}���\p>�o����� �Ⱥ5z~];ӏ�����.�+L{e-�#W�|��Hl���t!�����Ѫ[�Vώ��>c�=��}�A��H㋦�Y�sb���8�r9G܃�� /ӏ\��>���4.����%����؋��zG'ǆ%���
K-�ʮ|T0F
|�h��ΧSRa�KV%�*��%�?���?�~��Dg�B�Q���V�U�: 
���S@ �\z��#V�龟��ӽAT��vɌ4����lp-��B�F+���g@���A�iC��^��Ezx9�/خHh��  �G������+�ma�$� ��"�A����B�O�}e��i�inuMwVԺ�1mL�*�Ifk��ʶŮ���s�t�:�)�7�s�뺖�n�i��C���F�G�U��{�ʞG ��tz;vj�KJgԻ*��"�=��$��/�azc�]gҺ��g��k�&:�t���8��u3�c�7O~F=_}.��A<���o�=��5j�L��ŦX捦i�ыK���v������U�0���"�&!f��8�H�N��*�Xp�y�?�}04l\I�?K��0���X�V�Y+�T_&!99'�.ǈ��!�\�X�=s��� �� �پقJ���"Ury��I�G��f�u^Vulq�'��a�L�]>��0,�ķ����l6��e� �xЩ'����A���!V3w%��>���� ^�|:W���?A���;�����~�ܬ��~�u�u4��w_��Z��s��7���a�1�:��0� ��=L�B%+��R����Jojn�eO����Ao���p�='����(�\�#��G
YG�����o�J����������=����Su��c����I���i:��|��Q��Ҡ�\��-³h�����U�4qFAb�}���7�U�%A�?n[L�N��������w`��� �n��WD���zC[ӳp�q��y�|��|�9nh��[\E��P	,��R���3/'�w�=q�}��q�'��]4{��6�/�@#�ײ~� o��ߣ����܌�������Fޙ]=�����(�7W? Pw�`bid���T�+D�?u0r}~~��Y�G�h�Gj6��� x���� ���:Omz���Y��zOB�.��2;������;y���Z�鞏����؝+��@o(jY���6�hm�5Iͽ%���rD�\�4�6ּ ��wa�*SY扬Z�r�'�V<)�7���tyao�h��y�³O�hȆiR�r�(~� ��:i��������m�j�O�/J�S�ީ�/���-w����,�3#�5�_������н��u1uE��XҲMk9�9�yxL&��6[>�n��նj�"ƛȒ��zq����to��
��!h,�O��kt��n8��t�b6�)=���o9��MV��ӭ��$��|Ɨ��k���k=!�cO��ٮ�~���vךּgKֺ+��A�:����_a��F���i���ڌ#�0���\�|uB�WKW0���=���_w�ۦ��ӷ-ɬi:�5� iT���$S�L���ENԖ Dե�XlB�q߽�aͱ�������hu��oO�!��Yrk0���-{5iadx%<p6�ݼ�@5� i��{���Rί�S���=ӝg�.���J��:��}Wг��ҝ�]/[��MCɇ�.dt�SR��K�Z槦��uM��%�lWנ��%e>Z�Zs��S�L�A=R�Xw�rp/��[_�ͷ�_7�i={d�ZccL��/��w���>XL��E�o
+�g��_Su�c��� e��p���z5�>�~�ݥ��Ԛ?d�����I�߻sl��{��'�.w[a�&PŽq��s-=�ړl�j��P�����XY4͕{qC5��{|Q���f�U ��$����<a���r��ӪA>��6�>�6���KXL����x�%�y�n�/��Pݡ���e��x��������;[�F���/�����7��]��� ���cky��F��S�u{K??�23�m2٘��E��bfGLt][���GV��{��vm߱5�j�O�.�hV�V��C�u��H�0׵܋e�7������'��K�tmͦ�d���-���+e��3���[���,M#g���~��:��{����;S�}����]����=޷~:�X�Qa[P���L}7#W���/ƒi#"�L����<tk�[�z�Sm�SnWѮӲu+��j�%Iet���V<�JĠEFc�� _��њ�=��uz���ٍ������������=�R$�2}�� �5�:����<�t���g��|DԴ��n��t^F��w�F�V��Y���h,�VYx�<����.=yܟ=�:��M����V����k�r8�x�,
�w)%YU�)S��rh��S�dW�_H�DW�5KZwR����'#�<����s���:7�{Q������]W�_�gRdC���1����^4��еl�;5����O5iMKI֯��y�=���M��f���k�[��$3«!5�9|��c�^�H�چa$ʪ���l�z�C,��:��ҝZ�Z��b��ڴd	!��Ia`�Zy#0�*��ѐ}�������[����t.��Z�Kk�WGvK�-�x�=E\����k��j���LA��!1!��j��J�S���Ց/%zp$f+�f̕�Hޥ�؊�D��������$�?U:߳u��i���$�i����?~���i?/�8���G��}����j���}k��q�mOW�:�����^��=�wT�����2�l7�Ɍ?)<D���`fUi�����mS��׵j1�V��*I�AF�2�s����߂;���9׭t;��S�����m�?R�Ū��'�4�*��/*��AE_��e�o]��'�k����/w�սo�� ݧMfv�M��-�Z�Y��l�\��[�D�211���kQ��+��ʖ=�n�
�����f�]7g��knM����=>K5�*DYg��bj�G3��Kx�!XfI��3������Q���ܫ$I��k3H�J��7Y�Č	��'s3�{h�;���f�Y���?q��ڍ,?EvWI�N/Bj�x�-t�&]k�a�,�����32�l�X����+�o{�-N��{V��L6H��?����O�sn�1r>��&A�K����߉�u��th�ŃR�����Y�"*�]�p{P�,�<�\��^ٻ��;�=��5�w;�>�{I�Z֘��>��i���;+G�t,�+M�����Aqr�� #O��Θ/��w�Wv?H������5e38�SD��t2XwT���JJ�&`��F�j���Wݚ��ӵá��ҴpW��j�ԏ�� *A,��4�H�+��ȼ���I���l.��';_�o�z+�^��SP�ְ/�g�G7G��<Z2b�['
�^,��0�rW���:������@�kͦj$��	!�c`9b���(�D}�Sr	ώ�|;n�o��4�w�6�K^�{5�)���}�c1�R�k#F��G�G��s=a�]{�i:�Ij>�;{�wh���OE�9�׵��uuz�X��0��w����Kj������x�_,�+Φ��}im�.��Z^��}r7=���^��s������Y���Z��Pi�&�U�ت������czQ� �}#��@$���Z�?|z�ۖgS�{�u��uD:/�z������u��M؊�O�v�Q���v���B1����a��-��`�IfKQ�O$!Q�/١����<s�:7�Bų�ލ���1
XH{׃�'w�����h�_`?������|龽��>��oA������&?s5E����M�
�� ����i�3����zu&Zc6-t�"��V�y�bG]f�y#-#��_9�5�Q�v�y,��/�r�e�H#e��W��ǑP��G�<�r��Ǫz��5���MY�����:�Ru}�-_V�p[�Vu���J�MBF3A(JRUE�fg!��B�� =   ?   �g��z��� S�'����<�ET~d�7݆���ϯ���� 9�I?\��/�����6�r]���� ��������l�'����gƌZ��X4��A?�0�&��-�|� ����� [���9������E*n�x�� v
���� ϯ�y���_����5Y�;+ R[�ĝʁ� ;� ��}|�������� _������{"���Et:Ϣ;{��.�4Q�}���������F.��j=+�jy�f&Vd��)0�8�P���4���m.���췬m�[�t��01ƨ��"�ӼqKac�D��Vp����3�7~��aI5{»��b�yH��Y$H��C���U���������ѻk�/������t�Q��9v�G�t�l������ҵ�u.*�o[a��4y�� �������]oh��S�@�W��u(����a�K���實�I��l�ye�q��*��Q����c_޶>GBӼ���׶(@ �4�8bY/d�d��X�y!>[����^ܻw��v;�z_������K��>��C��M��;CQ�zw�-[�|����caY.���f2L}jzF�;R�1�5�Uy+��X���	���#7���j�:�QwM����L�#��i���:�*3z�<�d��H�-�O�=���m����^�����Kͯu^��L��������誅�<Vx�ҀDY���Z��Zɷ~s4��p#��(�^(�zH�_ВI�4�6��YjP�Afs�<���F%�Ϸ�B���x ��7gN�L,�]'0�YX5c9�r�%���L[2[Oő��!`��M�+��^��I�i����X֑�S3Q3���\|d���~�� �F��f�CqOLgX�/L���$id�||j74�"��3�O��a���>Y�J���e�Z-x���	�INa���Ы3���Jn۝��2XA%t{mJ;�*�&�u"���K)U���wc����2�г�ͱ��qU�zL�V~0~�0p8��<���7�~8*��|i����4S@h�B����cú҉�i���� �@#�W�V���� `��p�7�����ߔ�M�-(^dmF���7eQyP�;�c��F0�39vwY[(ɹ���fA���J��a)��zcY,�UKI�'KPͪ�vzSż�	�Z�Dщ	���Y�fy��@�Aд��i�:-�U�o�/&���ۯ�0YY���R�M��?ѷ��sc�7�P�G��<��c�5��Ք|�^�|R��9.1,�2Uj��]��G0Q�so9h�L�LY�$v�J�dI�YX�)�Rw����*���	�9"�y^�(�2℣x�ŀ��>��1��ڳ�4���ι%٫w�;�4-e���� S�q��-ՁJ<�͘v`S�9,�M��&�G	��=1�"V�1�5����W�/8䜂Q� d� ��,`]�"�b0�2d��ҡ&�Sb�&�
*�>���}1�_����A�p$A� �#]�����T��b��p �(^M����S���K�s`�
�"�
VoËS0���^,Ƃi��d#��@Pl��0�r�u[c��YWUdP_'̄"�ٔG����ٌB�3p2VB3Io;5Q�R{�c0�����du>��R.e&ID��.�Yӄ�����Ź�0ے�(æ助�~�B���]��<�x��#uH�;��T�o9x�BM|5�#�U>׋o0b�v)���?oL`Y7H���Dώ��I���͆՛�������0c$�x�M��D�5�uP�SO����$w
�A�nB1%<��&2��u���9�@o�E��}�"�&�,�L�z�Ҹ��i+L�5�3E�4�<��&�<�,�eD�#;6U7J�7��e|��.A���;��;( 1��^y+ff����*�j�Kx�	D��f��*ܶc%���q��aAi���J#��:1{n��7F � �G�1�,�����,�	����m�k����6䭰ܳ���A!�l��w�])e��4`$��+�T��$��`�<S��)@�U�&����B��
��y) Laը��d���#\yЀ�j��<�^B[���F���YyB�$��\�Wɫ�v���@�ǔՙ�p$��oL`�dF�H��Y�ysf(���
�	T6��T���I1�).���0�.y�λ�1�T)�����I�|Q)��u�4��cX��
����eU$;q2bF�B�L` �C�*��%GEǪ��|h���`�n�y%���`-�y-�ѩ
��KK%J��fFr�d�JX�w?�>�Ɵ(c3'Ld��S)��V!qה�!^@���vU*���)k'*�VX)%��e�
�
��c�dQ�K7n%�xC4��%�2� �>>
��\*�W��q�v\Ldn/*�^,#
eP�-6^U��+��Fs�M�^C�ٌq�J�,*�8��"�vE�($�7�Db~J��%�1��O��R�./�]R���YX�h��� ��ԉ�rvc&	,���6�e���6L��P#U�g�Kn۷&,�\𜇇�9�Ş��m�p`�c��o�8*�
��wb��i	��2Yw�p�S��8I͘�yX��� �* j���	VZզT�À8�<��8,Oʆ�V2
I�|���:c�J��(ȭO/�Wy�Q֟3�'oLd��1r�YqËi6�y��
�B�������c8Ug#��0�-Y�@!�����۳)�u㷦1ʯʜ��`�~U�s�Td�h�����/�0m�r(�G�J^G�2�xi���dP9}a��*��́=��X�W�Ɣ¬��~x~��Z����@y�p�ܰbۆ2�ig8ŀQ��Dp�7�lY�sja��B̚ B�,x�2+�-4iS^r��;ڻt����)���(�b��o��C�Zv^=0h���E���%Z7A��*�8m�(�����3Y�ϳ�V-]��$��ˏ���e��`Z�K��sh��I��~��h����<L��L�l��l�7
�f�lG��.��XyJ2q��g��3��vC��c'�c~.=�g�X�X�a:� J��~l�f��WcE݌�<~���Օr D#B�ڭ�:xhP�ODSY�]��| ;�ބ#�p	x#�G�v}{	�}�}��4~��u���CA���N��d�ONi�'Yɮ����D��&�戓�Q��P��������4J�#��c�g`Y�>H'f@>���ȓwt�E���Oo��[��	dBjؑG��R�@{^�q��H'#��Ӵ]��rrN��u�Ń�af e�4���Ř�!Vn���&7[[q���&�ؚ�ۏKP�Y��_���YIx�~��eG��\����ꆋi��t�Y�Z<��m�cy�~^O�	�����A�c��n��uL�����})�uN��JK5��-Zt\U��D`$���_l�-���Q�ph4�\�́lE�����k�����?����ͭ���6�^mR�{A��y�8�����U�(�z(��Yzc��[��������J��~��cF�д~�h��N���,��p��gc0�yS&���30�J���̯��d�u]a��Yk3�&��d��U��١���8�I��d!A���h[�T��N�zn��r�W"	���Z2w�c�T3/�ӓD;�J�}�����ptƣ�'_�Ic�N�0u��'�G�r�Q��z�kה+�O*onm�Y}s� @���;�^�P:��V��I�Y��~#i)��
��9$�8(�r;3�7~vN�����i��*c�?!A9S#p��Xe�q�)����t;	�iuΫ�m7����=��K�:�z>�}Z��u7�>f�z/R����u�o��8�$YM]���}��w�_�a�Ϧ�ܚ�	n,q*�(�$��)$���Z�=�À�)�w�M�z/+mm?Y�ކ���9�E>��	P�O�����:Cڏ|�_�g����Gys�n���Y�'����6���<cB�}OU��� Nuq䉏9B�okN[=��������7v�X���Mc,�B���ɍO��ċ-t$�;�H#V`{;�B�+�6�Y��=���+ojS���O�+�����	� PFY;ȏ�{[3��z����4{`������k�|�:_����n>�]O��Υ���/�jT�T����ٗ8����.=n���g�M'T�=�zL҅6�O�k��I5X;IXd@&��F�,�O.�k�Gj��ҵZڹ�Z�1)E]h��|(#����c��p�����)�[�vg��Ct�[������9��I>�Һ_������&Fj�V>f����⚚d�G��1ӟ�˻��v��5��Q��K�Zj�i:��Hg�J!��5e������9�O��ڽ5�����O�SKwO�.�(������؂&C=n�B��;��^s��/��{���������:�X��_U�����ug��7n�[H�԰�u=s��*�CP��|��{e��/=�YL�~��N�i{sQ�Bҡ���^w�X!�<��q|�v�d���a{��}��7�z�իۛM�[�bΑ-�Xd�W�M$k,�Vȝ�+���=�{�������d����/a����{��}9�i�s�}�wSW�~���N���gL�aU�ѧ�>��2�{-�M�8-�^�uGA��E�fZ,#T��|���o<gƬ�L�V�E'h�q �],�=+���wu}r�K�|R]J�E\"�$�w��%N\̎ݮ8_����O�?j;��ޝ�� n}��Ri����V�GE꾛��2c���}�����Em&��q�e�^8�J������]G��h��G��4����@�}�R`���$z�L��-�0n�C������{����-Qe}>�1i� ����,@T���n)Dt*\���H��W�	��k��a��O����fGI�Ή��ݭ�=̝q4���w���	�=�|�ĚdN)jL
	�S�z~���<]R��FZ6"M^���If�L�E;+�*�c}�7�߻f͍F�ҭ�H,[�1�/�[�g<��aX���PI��H_z�I�~O��F.�q�c����t��m���'���A,Q�c��H�bu���};��_��A��c]��h6ߦ5�۷2�=UV1�3F)�"��d�",l��Y�t�t
]�t�F49�{�n������ ��ck������m#��y�ʅ�er�?9~��4q�B�,��@��Lv��� ���jP�t;o �|���RQG�~�~G>� C�{�r9�0�N�"�8ǀ����~����������x����{ꚎL��cK+Y5����fe|ufi�*���m�{lQ��I�/d��1RT�Gz0#���=�N|��nҫ#A'de���R����G�ό��OC�7_�&����]Cm[�qtU�4��=It��0���|'IHЇ-��	
�=�F�蕌S]��Xyyy8(��y<(r)���3)���nX��BX���
�B pUy�A�C{�r����]���t�C��~�~�Ƕ��u���fS<�!�<<���8��T�;������ޱ��nZ���1�ʑ�^A��ϑ� � �O p�̺}:�Um:-I-�g�T2w�c�B� z෾O<ặLְ��t.���W����cc�ӵLigWN��UƝ��`����W/�2(_R���N��jK�V��c$X�3�gƳ��Gv 9R�ܫ��p�w>��z�i=h�G4q?s,=��А}�`��W����k��j���Yڎ���Y�cjV���=�H����у�5�[V��@f�,��%��i���]��YZhcT�x2�r�����?|y�1k��{*M~xl��Tv~��a�YT{�}9���6��gW�A�>��O�]����Բ:o��c3[՝�l0�?3\�F���t惇��j9Z�^�����{��8���v.�f�zޛ�M�$Bo<��,E�Qf��� ��I	��>4�b�e��jAL�|u�a�A ��0����Ҳ�������}���}���;�~�����6���h]1.��N�t�L12���>�k�W��n��%I�U�KHƙ�]�t�N%�@�vѶ4��Dӡ+�H��1WD��h�a�H��{�-Y�iڎ�TO��،,���K,{Xswt3/k#`�_]�0ᆺ�{a�}�`c{����p:�?�4n�{���[��滇����^ӻ���k�q�t�h:�-�^�����pz��
R����j���!�J�-�k��jt+��bf��-��xLWY#s,ȕ��;T���7�W'��-��h����?5��4�W�O#����$|�C����e�]�����/��L��M�z��:�G��^�ЛD��Zf�&F9����~5���9q���͐�7rA��_E�u����eI�)$K1���lJ��ӎ�&US�^Cq,�kL5�6�if�YU���Al��$���Hة�}�W�K�����:��n��1t��t�t�Le�XOP��Vh��V��X��/��*k��[�=>���o[�h�.�� ���
x�@ �����)6����ZUcG17 ���=�!��؟G�si;I�w���h�m�;�p��a�O�FgH��3��_�1��L_�>��r;eܼ})��ٝG6w�N�ۜ�oUӲZ�v�ت�}��{Z��w��w�����MEkI4ේ��+�Ϣ[h���D��#�e��o�w���4Q߾���{�V�G�V��>}5�f\@�b�2%��%�Y(=����=�ӻ��뱞�5ؾ��΍�Qi��{�ج�����fJb�uWN���~��:'Ma�GN��\��4��ѡ��<��E���A��F$�4�v���&T�]��Ƴ�:�D-R�[l+5�e�����i3p�T5�^������-Ŷ|Ve���ة{R�!��5��y�)�&h��&x�9�{g��J��.������{G�j�_Gu�Tv�5��l^�yuWto[`ZiM,��1�U���P��#������Ɲ��e���n[n�	 ����֔ bc;$.x��*r[��o����I�؂�H���$Vg4�e�U�|*2}�P�����}��m�z���^�4Z������������:�^��q=�/��ٝ����}0�Z�~t\n���J��[I�8��Ÿ���%��N7�ӭ����ح��t<���h����a����4��:4�ؤ#�ۉkZrV̊�&sstm}"��ܵ,���/��|�X�Mj�� S=-�m]J�Zb�*Z�%։��үo�������g�/n�ս�� �V�[���T��.�VnE��'Zꥲ5���S�%�!j�zrZ�r�1g��0���Y�^�ܔ��ޝ_�QR��PV�ky�{�4"�!��ı�8U�+r!�!i#��ZF��6ސv�m>�հ^T�6Yg��*�wRv��2I-j��dHԮ���H� �r��fk��5���gԟ�=����{k�؅�֯�oљ]M�u-���Гr/����9�p_%��^���u{:eݱ�S��2�}-d�#yJ�|á���yl�3�ܙ� �wN����دn+�m���I��c|�b��O�L�̂��	Go%G=�e���� l����%�-G�?���]3���枽K�����Ta�\�x���Ƈ�y��[���+���k����:��[��͠�c�K�1-x�/���W����xT} ��7�T�D>��7ލ����wH�x�-E��щS�ǌ2y�_/��� sG��]-��Oq�{�������Ov�����t�Pu���z����N���p�ɉD����S�60�;N���:߻OumݫԽ:��~��a�ZTh�H�N��ZD�X�}�4Ζ�Gcn����ޛ��t�6��+�V7CxEV_�T��Y�)�s�#�%����u�o�>���h'�E��N��b��X���Q�p޽Q�kzv��L����hW�܎^"��_O�	:���ץo9!��Ym�����m�\�Ȉ�]ex����%K0K`:2'b!��=�ғ��_QŸ��M�5�$��]Gt��2��e�5���sۓ=�f�_'��;5��O�oy���W[�+��w��^�ҫ�j�VQR�����ƍ��r��r��*���To��-S���iL�x��[2$���,e�4�k#S�`3R�!e����hMoW�SI�#�V
P��f{�����x��j]�c����3�N��GU�Fu7U;M����-�f)Z:V&�+��nT�;�,���D��T�����>����+Ă�Ƴ�"I ���X�����W_��Κ���꒱���؟�I<����=�S��O9�>��%���]��F@{��{�}��]S��������;�4=k3I}e����T㑬�OM�>.U%�i�º��+����껓M�6����(�ΰYG��I��+/�VH�Z��;�:�{�M�θ���z~��KWU����F,����f��5r�r�0��	<&F��j��%������^���[��� ꮙ��ӧ{{l��9���@���ef��1�J���U-,u��ԭ�-��:woKշ���]�4�,�2���b�}�$h$�̱ �#@B���ݹt��E�Q��N�X�:���^E�%�rx{PL�xD��(U,�C6j&��b��^�̎����q���4� U�oIi�\4\ly��Z�����|��u�Sj�O��O��-��wmMjU��W�W�.J�'s"��;bo��Mk᧩�Q�R�q�Y��#���*F$��hn�X�)�ޛ4_�������_�^��.WY�;��K��ҙ8�vWo���x�M���^���,/0uzd=sr�b���|j>o�(�V����ԛ:��vmOD��^Z����4�Oy�A'�ep�}H#e'���ޫ�zm���n�Tu����,�:�"W��c�B�@�BY$�;��}�?Q�h��Ww�O�zΝ�����k�Wǵ����]����m`����X���U�iL�Dk#^��4j�S�FHk�W�U�v�2�O���ףm���ْ�����-)�r�$����#����[I���r]��'L�׷ǢzK�S?Nꞽ����}�Ӛ�m4�L.����Ӛ����Ǟ�������rW"�|OR�j��jڒ;^���i�x��#��*|螹�e��y�I!nJr
�/���K?�b~ ���9�n��ѽ��a��h��o{Q�~~W��Q^z�x{������ږ���: �#���9�n�_Tȭ/��xj}i!�k�<�;H�Q o�#��<v)��Y%iI�A<�"BJ���<�����W�%Cf���a#<y��qL|Xc�Z�'��7p� 3>o����}� O�� ��Ϯ���9&��`X��Rv��ɿ����~���<� ��� \y�Yq$��n!?��%���̀����s�� _����K38�)�a��-�@���>�>��������G clV�X���l8���@⾿>�{���p��j^<F�&)�=2�E"��|�r~���	����G )@ֿ��@�C���� �~�� ����盻�sطz��^��G��Nw��S�گL/K�p��O7/��p��^���[��Խ����y�ij�<1�)�Zf_�>�=���ڔ6�ޣܻ�vuz�j)�g[���8�M�H���y`C��U�/2�{�w�Tm��m����<�j��E��4�bx���X�VF �Ѥ=�v;ؗMa��0�K��խc�����?��toGj0��p�c�=6���8�0����Y�Y��2n���ܚaٛF��7ۨI�I��X��IoT��<�'rduf�n�
r4�Zm}�b���e�rn�rQ��EHL��#�Yw�Pʋ�)
�¯�ww����v[��Z�Gi8�y�Wu1X��nC�#�����U�i�2el�+�v�c��xsn�#O��� Sd�k@:�򬾻[��cr>i������{J�wB�u]*��X��L��I�����$��p�Bk�� �k�/+z;�3�<<*d52q/��c�'���� �D�C1����NK�H ��	$�'�bI'�$�I$�$�d�d�>�H   �����@@@z�s:��G�Q-!$f��V��a����_���P_���c���iR�e_�gB;M�� ��Җ:S�֮�f�Rɨ��4gƽc�&��ҩd�+�����SJ�><��Y4��j�`,rg�)�M��f��D-!=�� zZj�n�JfVsL�	L�ܗ��˲A��JG��~a���f!�'r(X̩��^�Jd?:�nB/�6�*ڵ��;��/ ��J�*�fV3�c�",l��f�'�p�0*����珻��ne�Q��ɌvZ�$�o���-/���7��m���d\̿ Xٌ~CI^rQ�q)�bH�4M�&�-I�عP[e*��,ed#��:	��U�t�A_�t��U�آ��\y��+�Ȉ���9H����ޏ��\��l6c*.��gE��uk!��Z�@#����6q�ѕз���[�"�.�UN�]��)U�Q� �<�o0�b���Ƅ�Uj㨚�ɺ���t� �� �La&nG��Y�UcyΛM<si΍��bH,��䳩�����NBM�d�%y%'J9��b�&Km��W���c��c@1�U�|B��`Q��m��f�<@�����?�V��]�R�Tpμm�q���;��H�0ccE�5x
���%KLy1��h>�i��Ȯ�p�,��[y�)���9��T�����a4峾��y�}1�QJBTU�Ѕm}�MEW�-�,&�Uy��?,�є�U��	��x����[�(8����c%���+�/�"�qӔ�>#��ܯ-�'��~}1��l�-�7����D<�6�Ni6�_�T+�~�0ه�0����B� �67*�n�ɑ�A���G3�r���0�r���9jX���49U�9N��rN\@�]�1��Y�s�Y�X��Zb�5��4b]JY�eB�k�S`�����)�C��(�L8�]iaDA�2[z��b��ጊ�8�6���5�������.� n�Ǌ�S��2�abhǑ�d;�^�2i��l�v`q��x��a�	�ő;4ڎ߱�$�g�IyT���|7?_P@B�jY�3k?�*��&�����6UR�8n �|�K�cZ	��J�_���y��ҞO����2$�RHf0g ���Hގ� �� �"��*�b<rķ'��!��y7��=)�M�if�(IyՁ+�@� C���0�YMҩH�5d��[��O ��d�\
UHR۹oLa.�^<�ʮ�H�B�$���k5Ln�Q��3o��X�B4x�O-���� �U/?@Q0��vNc�8�%��zα���ζ�
Jl�#֜Z�W��n�f]��Ɍi�0��f)Y�SV7��`|f�c�HP�8��n#��3v�
��P����eQ�#P>�g`�*w,cF2y(����"�)l���ʂt��φ�鲲���cʒ������כ�ٚ�km���  �K͉@����WD�B��l:PJ�
S�HE�e�[}�cI��FQ��U���\���ug%&7�U�$�Ō"N���P[{���u����g �j�Fc��<���!�yS�	���y�PV\W����^k�۟�Xm錎���$�G�[mV�(P�ɛɳ�қnC*;��n�)��#������7����FI���Q�0ݕ�|x����͈CLW�W���(��YXn5��g��I��ĩ���rO�+�MTvW��ԙ�T*����MW�@c���a�X3�2Y� �<�� �U�(Ux�����֮:���i
�Ʉ�QFJ�HY �4;���1��;sWFȣ�.ƾ4���ļE<錠�^A`	� ��pA��(f��,gTdJ�-)d�h/�����er�B/�0��&�VL��j�P�ʄmȲ*'u�f�}1�3�K�ZygCJs�Ȫ�N�&� rg6PS�V06��Ut�	:	�F�,�l��J�<1@!o��
��X�Bk15�o�zX���f����e�KH���8���<�RJ�����F�-���f�]����:l�Lec/Llu8��5T<W����~;���u,�1�M�b@��j�-I�@⟷+*P/><�7
�fSva����mi��T�C!JP5&�z�J�ړ�%�٘n�qOLe�y.���	�Uh���mWC5��aUܱ䡸;	,`�	G��L�\�8���1:��+�r�q;6e#v2�Zdq�Ȅ/�\:=q�VQRh2���Ⱦ0���c��Z�e��s�bS ��$ZK7��@��������1�����,W�f*����C&�i�!�H���AdB��Lrx��-L��c4o���'լ��c�'<W��N��j���m���R�wY�����{P����gi0Z�&u!;��dZ����i6��  Ϛ��Լ�]lf�*u?@f�q�������q,\�'�-
d�iVmЏ�F_Lg�������15M�5n��Ҳ�������蔎DS)YO�&I(�5fF! �iZ���݋Q�/I�݄�D��20��F��x�V��!����N��җM�(C�П��΂H�)��2# �ȅd��de �c�[}sZ��^��������l];M�1�V�&`�(���hNZ~��&2x�P�R{3�Ogk{?P�`}u�Լ��c���;�wIAٽ�)z������f��wMڌ�m.4*�&p��t?��s���� ��P8�ˀ|}��Q5l��tFp�P��=q���;P���}?U��rt�Th��,�z`:S�rPJ��-uCq�v�;Q�=j�*�����E,����b����"��ݻ��{��y�����K �yY��}2�f��@;f�T^�9��k}�vc�z�Wթ��m;����&����]&�m�����f��畫i,%�!�"x�g��ѝ�42n����դ�A-���W���=�8�1�lh��~�Y�s���n��ޚ��\\�M�e�`���d��0{A/T�s'?Jȣ��}ؿj���.����>���\랼n�螠�ms�H�-���h�����C��t�@�U1m����V��� ��������m7K����`��(��j֡=i-��'��HC;����2�i:?�������=�n�~��E��tGv
�+N�
�j�Z�x�b��4`.S�ٱG`�?�g����~���}�w�tZ�M�7��,<q��j�~��i���鉘3�
15��h�I�sR���c��|nM'�MN�:-]�i���v��֕��o$����'ҝ� G���7��
�I�-�T�5��W4�+�ݩaH�C��,Y��IWj� ��L�����������:��;��ӯ��Q��m�|^�W��J���K���\0�����sf�\��nG�/�M>��M�T�M��*L�0{f��Xk�JS��H%����U�M��mZ:��ˡ,���i��#�W��UB��G��xӁ��{��]��'a��vS���z{�Z����c'JкW�t�;Z�v���i�f����>7��ڦd�<g����8�C)�]>&�oO���b6.�MS�����VEEe'�
����6�!!�RN��9����ַ_��W����u��Y�����fD�+�"�J!O<y�d����u�����0��Ov��[ӵ��zWQ�_�:��4�E[S���)��:��</��L�w�|����K:��7.�] Y(���kޥy�@��5�)��ya$�c���6穽%ۛgB�I}���=+��Vx�w�1�"��e���{Fh�X{��=�����{нO����Pf���'����.�w~��n�l�7JR����d�ĝE�8��e���
}[���֫_^ի��jOKf��V�>�����Q�"C!f��7�z�o��J��m��>�7�t���x���M�����G ��TvX����?���^�}��V�ގ��%��ϤTv���[�=OQ��鐸��5�SY�W��(NU�p��l��
�`�o�-��ts�Qɲ.O�ŬJ�j�qL&��)��U� ��ڨ� I ���]Z�ȷ���kK�94�� �hI~�2'|QI3G"Z.Y����i퟼���=�hݟ��h��=����Һ�����v���&���Э�2r1�Qk.E2��r��ŖK�-�խ���X�����a�&�n��d�^E�~��ؔ���,�)=]�}?��6��np�H��]F9�˪oT��0�±G$`��$mg���kݭ����+�qz���1�>�W��W����L��������~��SQ��Z�E`:va��U�I_&X���b����յA�n�	<b����URUd�~&+P�}ʷ���!�iuy�ߴ��:j\���Y�R�+$H)��3Zs�#W����sFYc���H��Pk�}35e�L(���o|��V,�����@ ��Ֆ��S��O��� ��珷�s�̖�~W�H��yq�����8_�^�������=��O.���|�0��fu �W00��)��g%~������~MV��,G�-$�Y���}�?W��<z̧N�i�NyuX�eIUP����q����~����gt��Z�����.��=+K����V����p�a�i���i�2�p�_B�/*}h�]�]����W��C7��(�X'����n��YYx璥{��t-M&��	��
�Bd���)OkGa�/�YHe��r1zgQ�VdOA�X�v�t���k��j��Wo�yX����g��ꇤ�<��UM�y�u6�ۻ�a�� c����Ȳ��$9X�����4�A�O�8��cn���R5*NC#�<e��(���-�������y�n��>��vӥt_�0�Nn��A�չ�TE�n���R��xHdд����|����=O�����O#��%�8cWu���,>��',�y-=�OQ�����"�O
L�B���<�8'�Fl����k���Ϳt�;����v��:���=��u�[��ڮɤ?.]'�k�!�7]w��H�>��2uJ.��{�Թ��{��}����k75ہWJ���-�{��V��=����gܭV�qj�&����e<�.X �����2��U��hY�W�����d��zˬ��v�O�g����^��]�������'�o�N�Ң�_u}��K��X���~�̮?J�GQ�!������Ƙ���vm
��M�MoG�{�h6Ht�0�;�4{�L�F�@�Kʱv�/�/���^�j�ږ��:e�Z�݁�ڨ ���'�R��O���T�7�Rʽ>��}_��k�C��캂�;���?n�~���g��M��k��Q�gZΖ�+�ݽ\\�c
t���txx!Lb�����>���$ږ��>���:Ƨ5��a��$��2~�����1喢ܽ-��V���]�H��BIe�|��ؤ�H$z?��^X�8=���N�on�E܍�����.���zˠzK����и��<Ο���I�ދ���P�7F�>30�6�;gd>]�}Q��8�?���Y]>�ͱ�ڱ؟æ�n�rZ�*�VKW�i�Z��Cȱ��{!�����}�*ۙ�_ԬF${��_�M:J!a��|��ր/y�9y�(<�7$��gwc��w��c���⽩i��N���K�u=�}�v�����t�����y�*4���7�5s��v\���� N��=�0|Z���w=tڝD�i�i��6��b��XcMoJ5y-G#E$V!d���NDl��X�d�v����7���5oh��y�Ѵ!i�]:�[����F�I�3�ad&=��}��D���_�������u�:uOUu/E���>����������h�q�n���9��-5�=���q���L�m,l��Ű��;W[ժ쎠HZ
W.�]&�r�<z����XY�Z"!mQ1y�'B��^�Y�0Xֶ����C��i�I�}>�*{�Y��cI�W�jz�b�d��6��� ������7�w�n���պ�t|.�׺��� �}��5����LI��/ҝ5>�����%�5ïO�S�-�������c��]��K�{�eP�mt➅�^��� c��U�������jv�َ��9�W	YUN�t?��\غ.�^ר��Y�w�jR��:u��*ԑ~U�X<�<c晧g�2�f�����=����F{n��t���H`5�+[�>���տ��!�t�f���:WX�k�ٍӚƁ���xyzrx5I$ƒw��S����}`��v��Ь�aWT�r)u}�#�4�nf5%�a.ӽ�$��1�91� ^�m�콩�n��mq� ���H%-k��p�?Q����U~�� 0݊D������7]v�&�ҽ��#޿xu���>����o�=�S^��}6�� �� v:T:�;+�SǼt�cmo)m�Yi�eaKpv^ű�uMKJ��3j�̡e�}� ۭNՈ��C�uܡ�QR�Z"�+k��ZFӥ��[�U�Sp�o�������n{<�Ҵ�P��,�
�UVTB5���op���;:K�7���t�s���t'[�^��X����G�8���C�{_ڙ1^����t����N^f>�mW0�?���ҿ���zA�l픧r�0OZĢŘ�;�G�RԼ$�<�j�;
�J*�X��7�֣����-�W����:M�:�)�J�b����-"�������.�7Z�����u'�L��>��o;w]K�;���i���Iuǋ���^���|�.�\�m3��C�eS)�#��t�.��z�v��MEmV����b�z9|���vz���~���($���]FdZ2GdY�Ũ���q/1܆bL��7�2�w^���\����?��q�]�ֺw2�GD�]r�?���ˎi87X@�tuY	�Q�M���N]��]�	�U��BIuj	��+ܯ .C ;Ow<q���ޙW{��e�mi��
����qYdo˙�@/pbOks��r 9���+⾓������I�</�P&��'��|,X�2�v4znn�6Æ~>��}�Ψ1_RV��nq|{� _�4�gkƺލ5 �Dh���Si�Ft��j�����B���;��Ycf@��]�^}"�_-���"M-P�WUp�V�)׋����*d9�~�u� Տ�=eҾ��mc/ږ��u�op������-�`�<�=;�����0��e���V��%/�o��pu7Y�i��h��yIX��%�'<WJ��If,�L���t��n��.�K)i2�ۚ�/�D�`J�<��l�o��i���?c���`�k^�;��9]��/f~��������|-k�p�WU�>��l��X�V����������?�r9����}=��t���՝��vZ�ȚQr�U���x���^e�#U�)� 榷�w��kp��'�r��kY�3���ڈ7��$�.YP�awg�Q[�99���}����^�� ������k'�r��w3�zm�=7?���a^�Q�����ME�d�IG1&3�l�=8���.����ZW�VEc�&	��q4�����?��
��O_K����uåuwj��(� �jq�[H��,̌��4��AڌÞI+λ������ x}	�N�{��L� n=5�ϯw�u���_к���[W�=O��Ń}E�rg��@��l�8NM�]����u�u��>���v{5��4<��(�k���#嫲ԐD��C�V��ͻ�=X�{0^��[��`3Y?��8�yH�o R{��p����7����<_j�!�}o��`k�-�t��.�ǷTI$��U�k�X���Y��ҟ���FE�I��uS��O�~��P�
55y�Hff�(��|5Ex���Hx�"��>�؂���b�z���4�����ҡJ�Ȓq��Z��H�G��<ά�9-o�X�����/�����Йf��7���4Vд�=2��:��\��,�_&���L����N<m�D�:%�t�_Ӷf� ךJ��X�v�s��+Y;%�}�ڀ�~�-�ם7�z>��h�sn�倥I�T�Ko�X���+��O$�������r���~����_oڿX���ܞ��������Կ�v����T�N�����N�Ӵ:cbb\A��G��j2糧��iڅ�SS�>��u)dgy]�R9%=�$j�2���Pq��#rw�� ����h-K� T�8b�K_縷�!�I727������#ޟNi}o�}������;��oQ�gWh�N>�s�A���4�S�]Fz��O���2d%��Wek�al�姉V�����d�!��T`A �� x&!�a���Oҡ��UO�U�o��VrCF̲9V�3T}��Wٷf�����X�~��HghK��~�:�z�Gq5ZIs4���z�b��T�z�gS���f�h�������+�v�W�Yé�R#v�?F,ݜ2�%��F�*�'�r��Q�a��>9F�r��pȧ�<�~��Md`��H輥�=����zK��a������3|��tfw���)riOd�N{�w]����ws���_a@NUC#�@8@�?���� ��y>�	�wNd�R�B��m��nH����� >�y�~� �`~� ����3�6_�?U�Ň��;'��������������o���������3!����z0�w��#�;z��y��^���鲾�p��f@��A ��� ����z� _�^�ߣ�$�*�T4����`�� >����F|�c� \�t�Gu�r����w�Λ�:ӯ�˨4Ν���/#X�.��u{�LѴM75su+��sU��r@�ϫ�!Y��o�K7
;�����PX� }s��8�t�,1���Tw,�(�$rH߬���K�;ɪu,;�К�@j:P�:��{���i� ��[�r2q�˧4N�l���Kj��Zej58H��v�aX�V����Lc�{�|�1��~�CnW�^'U5��	uh#V���a���/���ѵ]kC�/K�)�֦����ϒ��;�n�x;�~��c�k���F��y�� Mi����1�13{���G/)�����=Uy�̰�ԭ/NK��|�Ww����֦�>�����^�nyc� }|}SK_Va�b��.��辵��In�Bݜ���O��QI=�C,M)#>Y}�~�����݁�ڷ.��]+Q���1���z&.B�����3�m{[F�c�Ҥ�b��:��nym�����i�y��[�[R��u�#���*x?�����V��ҵ�׵i�U�r'��;;#��ף��� ����`�ep�b\�t3kz���Z✙.&2c\�yީ�K*(�wR�.*�~�b��f�t�G�鉦<1��ى���!���.��B
S�(�_�}��z�h���>���}2q�uHb��f�Ɏ:���ea�uY3�yo�#%�8Z��KV3r:����ʪ{�曌l|��6�����I�k��Jf���Y�fWcjMьގ�v> 2��n�"-6�$���J���K�1Z�� |�pvDV3j�`�O��6����8;�f���h��	�~\�����<��˦��t��-ć�ܬ��r��y��~~̟��9�$��>�gu���dw�ԣ]��,�%��[/)��MK��݌���Uֻ�?���z��L�$�\ԑ��n���L4�_5&�����*�Y�"���4Et |� ���S��"̷d��Y2
&��`�N,�p6`ILc�^	)Е̽&v���0��x;�`���Ā�y1n�X�
��gfx�5?f�~*�6SP�ʊKp�eI'�F7�Ԡ����U|�E���Kc�ǐ��M��I�:d�cH�y��l�V5�V3Ui��<��O4TO� �<W��8
CUX��!\������iC��K����H��I9�!C5��~��IB��1¢��_0O!>��Hd:/�S�<~B��I%w����j@w�/� �XʰE���d���ɠ�U�ǰ#��(���� '������Q$��*����@P�Rl�f�G�<T�?��X���b#��4��ebѐ:F�8���T��!����Z��3f�2D�FH�4�N�X�	��l�/�2Y���Dw��&����#��9������}1����*�
� ��:��m�S�|�� -�����Lg��_*�^egH-P��	����	�bȢ�R����aM�,�v]�2��t�+mR~9v .�X���rۚ����'Nr6�%�͗���/�c�γ��ʵ2|S�.���d�f�,(΁��L�qa�f0�ƪ�x��:�W)���Q��F�Ҩb>��*|ﲏLax&��D���)8Y�K#JfSbuf�y $����4JKP�ÚN���l�,��7Ejp($�B�x�-�`�� �6�j�UQ(���ی����M�;�#e���<e��(>`F�R<��Vgp��m�
 V؝Ԃ��ьQ��*1UϚ�����9��m.k6Z�'b�\�Kzc+
��s�QJ:Wi��,Kȿ�@O� ����n7c�x��r��+�>U�d	w���ʋ��0����c�nlH##�[©��2���Mx�*!upY�Ō{��Q�6�5�1�H�UU9;������A��OLc�#��u�h�
R��M*��+��b�v�A6}�,�Ǵ�(G%��
Ar੒M8epD
�_��� �� ��8=�芊���U�Fqc��4�@i8�BX`�0�6_L`�*�D������@iO"2��I
�Ef%K��rZlaUV
8��⿑	�2��r�����m�"�6���2�M�Ŀ���h�P�z 9�ܦ�Bn�J|1�
 �E��*�� C�2˒X��"sۙ��I�n�=��dK��/*�+�Q7m��گ?#*�q�v��=	E�Bj�E����4V>^Vo.�vA�G��%��c(�vĚ�*�D�J:QL�Z�+����e��'bO-���L�;A��!4F�[!����%N��CәwUBN��:�Jm�iI-8U^AVj�nu
#Pm�߉q��ٌ ��x��U�c,���\�g�a�r��t�T ��D�%<hJ����
?�թ����Gr8�+�&,����r� r�M�y�,��؅O!@�+ɐrf1��&��ƎK-7�c9U���6�}��bN;5�6~ag*�"����f�n�~�� S�ޘǦ8!iG�3_�[7�ȇgZ��Ȧ����;�l6c	���s�N��
^�g�:�e�Q�R���'AD��8<ơY�d�&�QE��������0�[ġy'ę�����p���FlP����|tm��֔m�F�+��������j��Y���3��VO�V�x��)b�B�݌�	E�bD���:dd�j[�)<��$|�B�b�{�~,b�sGс �K"����w*�(���.�F�A�����TI�\�A�דs��JS���Y��U]�Wc� ?,�* ͣj�x�Wueq�����c#�=6I�vi��v���Ts��M���i�
�$f2'��fZ�Oo2�<�n����e�Zr���U��^&c,��(���-�K��rv	��f�N�� ���xlU�g�Ok$���7�x�|.i��@�r�T�3�4���wV2�M;��)�&Ӎކry�ԯ�V��y� �s�V!�1�;]��q��'�[R6\~YGj�!�nF��y����U�Lf�~��Tl��9�!�N�[%�])�@�Y�Q�dje*xg��oő��t��a-s3��sOV�?#9�H2�����;"鴔��o����}1���7gu�2���ic&@Ө����,�<��᤬��|s[��c5KP��mZQw��4�*�:7)��;4�w��eo��X����� {��u~.�ڞ�mC�ڮ��o:����g
��_��K�ېK�)�n��O��Q�k{rF�4�f>��f�)��wF'�M��b��ӥ{R�p鳶��uӱ5ʞI#��o��y��l}I��h�Ϣ�o� ��k}��įzK�1���#�<>��3�L>���NPh+�o�f��T�lI;!��t+4�I���T��+a#��~�.�c�|��{�(�Ӛ��morӚ�E�pM�Ye�j���Lg�̓	KK�L}���)��fS�Ϥo��j{U>���鞢�P���Z�K���:�L֚��Nf��hYRi���\��$����V���;G�:���dW&p�Rĳ�"C���]\ G2�h��@�N;mk]8۔u��Z0�ɴ��Ow�;��F²�N����$��\3u�����'k;[�}	А��/"=��M3�sz�3;Iֵ]�$�+#��N���T��*�b޼��I��,��4��m���K�`�J�����Y���o��wJ���EYO��L��EԷ{ɹ5�恪X�2ߕ������Z�ʆe�O�\�����~���z��%��3G��qe�������:NZ��V�]+ZǾ��};'�r��-����bΌ�}B���{���]*-׫\����Z���k�K%�������,�D���N��ӏ��Ϸ`��ٺ.��ߍ�mX��]㙠�w�1����H��^�1�Y�:?Fv#��n=�{i莿����B�t�vӥu�3�a�J��S]CW�Kg�7^L\l\�d�U�t�:ؠ�m��=w��j�����dU�jӹ��i�,o㍡i�^h����r�)`��	o���z)���lGGX���mC�ʔ���n����֐��ٕ����4Wws�l�?H&'J׮�����=��W�z��tf2���<M{R�8yU�UB2����1b
�?R���I�w��t:�R�8��3M#z-$q¯V$y{����f������%:pj�7T�)-%�c�W�#ؒ9��aF��r���.��?zK�������s��ͤ'Uk���m7A���t��7M�be?'ɇ�
b�b�~C�fE*����Hn������;�jg�<I=������z��=���N�70#��#(^��C��o�t.nx�ԧrh�H�^$�8�,s<0��B���ὶT�VA{��/�m_�^'���}`zY��Q�;+H�z�����#v����G%��t,��)0ZrE�ɯn�T�͸���؊z3��*yk!�Iwj�eX�NO$���N�-Y�jjڭ8���q[�fB�'t��	e�C��*��ܞ���:�I����s�Z����],:�VMk�r�q�-�_"�F_�Ue��%1�'5��t��`i��<�h�F���0�~������'O�/����ƈ�CJ� `�v����,����)���z�B�1�K�=��z�Z�m��몺h�91�j5����z�I�	_'Y�􎓩�)���^m���jc�������]�k@��&���S�V���*Ա�5)�!�h"�R�
��W<,NrO�
��~v���Ў��k��L�!pk��&���	O�2)�����_@������:�*޺6���N����Ԇ��ǝ���T�ӝxۅU]YF��Me��He��οO�����x<A�O��E
�����H
���%A �@b�9�zw�k.���s�3V�ǏQ�غ���I=?6|�#U����b�sO�������/t��e�.Q�����������0�Ǳ�:շ&���=Nk�U�G �q�q����s�ǺZWa��Lѻ��=z_QO�ӽ�c���Z$W^�u:٥����.� �ZE��f�N��;��`�-�y'�%
ѫ����s�s�w���i��?/&���G�k#�pyu��܄~��=�v�e��t5�}M؝����Y�c`�}ӹ�b�_Q\$N���8�UNmL���;?(&&.���{����V��iuV����c1e?�㷇�|,���C~��Rܗ�O>�_�jW�d��l@1��$�? GA�rxP~ٹ���|���S�����׬�I���i�~�i�^�� �7McE��3u���t�QOM�oa�yYs��^��s3��˴4� C#S���o�R3�[��o�sYy��Gk��|�[S��Gfc+��X�1ֵ}SiVm[[�Ƈ`vǧ��Ix,���}�`p��ܒ��L��/�d�?S~��>����=����S����}lN�v��'K�C;;+�]��5*�t�[�J��7�6�35��w¬qiq��}ɶ�5��ul^�w��eka[SM��ʫ-@*�RY9�8�k��*�c����47vV��.جT���gE%	)f$<U�v�4��R��	������k���or�ܬ����e�z?P�]'������˨�C�N�af���o�W�ӡ�,�kZ���2
1ԣ|S��rt��ϫ��Z�j�3��ۖ$��f�E'h+�ך�l���<��61�g��\��GA�uK�W��{SQ���Ȕ�j�,Q޷fZ� 1,p�4�0�!�]�^̽�B�QX�Ʃ��{��l��:��5�~�msZ�����gߏn���c�jz���������V�� ٔǶ���f7ˆ�s�ך� [�tãj��H��V��DRi��5�.c��ji<ѕ���s#�� f��2,��(Pډz}��Zۚ���I`�MR��I�}sM����/*�|�#��_��ڟvu�{]�ޅ�ߧ���}�����}��R���=7��н���=I�ùZ7�`���X��ߏg}C!c�y�p�t��i�M�zN����}Y7Ҷ(�Z;��㱭�Z���)��ޔ��<W7fB�G�/R4�m�-7]�v��Ц�O45X�.�դz�C��m4ZF�0��Լ�O�a�EC&l���ޞ��f���h=����.�wC�z�/ޮ���C6��Ϸ���ݝ�/)t-H�����Ա�q�%�(�*��
>����}8��I辠�����E^���,F5
u�.�����Mh�*�d��2��
I{��}u#�[�Q��G���֒��#Z���CQhU���L��d_�*�6��v���=�����+��틲�sێ��f��ޛ�_l���i}��2��4����S<M3��l��/K���Rư�X��Kֱ]������M�wF��/w��GG�lis7�K^��}=���e���K�f���R���L\��C�j�+K��U�F�ZwE�^o���Z*�s�#'9�=��	�=��ܯio{�Gهy+�h�Q�u�{��a�����}?W�w?�Z�M}��"��?SЙ:w/#�~f�*W����ѽ��ΚmN��=(��Z]��oH�jh5�i�<�F�F�ƞ���*ji%��e����4�r�+X�V��;o[;%ıڭ���C-I��	/� \��]ĥ�KJ񬧛6��9-�};���t�k�һ��]O��wG�MOx]O�5�=��t���V�~��Q�Zf����y��M3�[�<�WW��D�1��l���t˩;ߧ�N������mj�<��v�e�����tT�\�4�d�#F�ݝ��U���-��n�ot��+�Y���_����hkY!=��k��qL��c$e9��C�5�d����:��uڞ��ݎ��֯�wL��;����m�YP���Ӛ��H괾V&e�Q����"���h��m�j��uՐ�*�.��%�<Ac�\�R�c�v�h���I�����m��R�u(��S��t�mG!h�Rd�(y��V���X0`G�Fxo�+���ϸ�w+��^w�G��ө�˶}�y�L�c#O��2���� .�^��2���u�<�4�B�%G^>7mξt�X����V�m[P-;��F�N�!g��QŨB�c�w�H����y]����.��5��[m�w\��٭Fi"���h�e�b+��BM�H]�A�Ut���w�ݟu�CО���;��7��/�p:�z���-Jвu�M[[]!��H���]��<���w���z{��&��Z�NvF��nhh�j���u��8���!��0��������~���>��lm�oV[��bO�eP����J)-�����3����)��� ����i���O�>������iu��d�C��kd�[E4��i'�|����9i�_$�8�>�n��j:�G�[Ho�qؕ-�I0�a$i�V5�h�M'p�!(s�' &@ٿ����6i��"9j�F��j
�'X�O�H��g�������N}�tz7D���s>�{U��ߺ=��2��ڝG�0��js|��#)4,&�������ȟ6ʆ6�H�َ9i����˨u>WO�%�U�*O#,u�#�;
��؉�EȤ7aTX����Q�{
{6��V�+Y�	�"��"�3�]�HC �����w���s:�x�����uT�����]�����{����:WQw#T��kt"�+_L�d���_ʍ�dI�~��[B�K�i{����Ɏ��Tא���+"�l�!$��:����W����|o�U7��m� R�@�4��Mm�-ڑW2���B}`K'�7GޯY{������� Iޛ�Rt���y={� ��wG���������3K�L&��=GJx�u(�.>9�1B�N�_����i�e�[-�0S�P���DAb�fqZX@x���H�J��������gU�N �i�<ƭh�����BY�B���b r��3��o�=��'��n��C{o������5�oG��ӣ���B����ޜ�2)�+�D�S&
��&�e���g�7>��F5�%�i�4�؞X��4�m��<�$�R<.����Ĩ�$�z��ӫʛ^��bIc�$��8O*: %�хfC�
�Ǭ;��[J�ͮ������4��'Rat�NGH Ϙ���QƮ6���y�K4�!N� i[g�s,Ig}|��MVI�lw!�p�Y��4k�)Im��� ���;P�k�I\�B�����R�PxPv�L��s"���@W��O~���;י��v���߭?�tV��>���^���}�֥���\�C҉���[�N�j���F�޾������� )��d��֡�`��;y�c�{�Et�����CwU��B�������"9ѫXNʲ^3�"5vY�x8ā�#ۜտTn��}M��鎵���i�ڬU�޳�:��0�?�ޝ��YUԺ�X����I��<�v����(n�7�J[N��ڔ���<>yɛ��o%տx����2�?��&\�n+�v�ΰWF�A��L�����ʔ�B�O 9�I�_o^�=��~gW�3�t��m���4�\:��m:�(V8�m�\��t�9�ͼ2��J�B
��-&l���=#N��k��'1��=�YB%���A"��8�
yʺ���E�ժ���>�^$^8��ra�x>�Vo��j}Q7Wt_�}:�;��t�}=�a��SS͊�oc�7�B�Ƣ�Sd����J�Z�G�4��G6�*���t�L}��~Au���D���y>f�ב��O�J�Y�d/���x>��>{QG�����h� SuF���G��WTk���k9���umcP�Ե,�Yۏ�ge;=x#*/�TTUEEG���c���� �   ~� ?�z � PO�}��?�$�s�0`���a�;�6�A]����p���={��� _�����r%�s��[��`���� o� ��������矜��� �� X�W�.�(rWfS��>[ḟ�� �^�n?_�����,*w���ޟ]������� ��? � �}�����y%�S�����ɜ����#��?���_^��G���$������d���Ϋ́t�;;5)�+f&.K�cee͚ն<�N[*�$��Tc4 n2���5���E�v�Qj�Ff	x��,9��
rn��HUVc�Y��wM�zsꚤ���ZG�|���
 %��!�o���z;+E�7^��tlv��7�u��M7������,܎����WU�!��ˍ���c��'6��lF��v�K#��m	�nޢH��_X��W���ZRL\�~�l03��^���t���Y/k�ɢm�Lzw ؞2=Ii����N�*$`yd�w_�gi���_Bt6��^����I��im��r�*�Y��N7j��4�v�����y�C\�ŕ�A�f�O��Rܓ��BR��!#�IfOf� �M"���*�[Ji5$iR��i0wDڏbx#P;ZQqũ�'�@Mh�,���9����{��mO�z�q��u�Y�,KV��D��NJ�c�]9�NF]9�㻰�1&����s�,���OpZ[Z����$�W��DPD	�>���n^Ww%���h�v�U���xĭ�F=�X���%?T��'�E�#T@F�~�����V>G��?%�֕Ȅ���ʔv�Q�M0�����NK�ϗl�-#�'�1�J+��	���v�\HJs8�-C��k����:>2ԡ\v���ӥ�dȦfT�����Z��:��Y�H�l����J����1���؝��\<������Ӱ��Qt���+䶟���*��Ǣ�~�Z1��%�����$���|&�2E��d�����zVv�Ϋ��MB�yMّI?R�moL�^,�?�xq�)�a���5q#�����i�\��~�52~�2,f~�XU��W
Y�i���+�iy%�ƭ�lBN��Dȣ4��jzc2��1��+�ǝ0�ߺ<3�<j�·���v-����&��X�[��8�J3dU1�.��.c�j��>)? #�"�y����c.���5Ez<&�>+���?�b����Jc�v'�c��C<y+(%IX��@)�GƄ�^�N��o'ħ�22 ��V��C�.Ʈ¶�I�*?�+*��o���L�E���j��5�Dg�y)�v�eP���!K	*�%�V��O��!ك8>YQP��H!�X c$s�4UU��jՋ�F����.w$1�� ���(|��/Đ�6cI͟������1�n��%�W2�������_j��M�^|@ �}BHcEX�Zy��(�����Ɣ�*?m�()�eo"��0cZ��Bx�`ʉ��7��tN^E���7�"v1מC�,|�	�FoL�?�Qy~f<X�'bX������0Y)b�)cv{�4,��K[���0H�E�1��D3�,t��W*|�M��!d+�ƻ	�2q�I�wc��?�-f���t 3;Ju�Tf��(IPO�LcYf��͋0�V�T�/3J,ځ(�W��K�6'��c�GV*�B�Hc�i'��~ٿ����� Ǧ3�>'�]
DP�V	5jD�*E�x�л*�ԅ�`�+��h��v��R��R(cBL3�
7��~\1�Q7�W5��ݿ#6f*7ڗ��'G�)_�� ���`�)I���tI�<x���m� �گ� >KQw�X�$b�\d�M@iP��Q�Y�Lm��A��r��c��2}�M� F���Ӗ�6ɩ��G"^���� �����&�|�v�=�-gǊcԞ'�)f)�8N\�c%<E$j����AEy(d�;+��%,|{+1P����%�Z���b�yn�TtS�s<�]�Yl��e**��c9eҳF�*Τ�����\v*2��NJ�_e
M��e��g�Ȧ3�/�p?�S%��.���ۈ,>��X��vr�b��+���j�(���9Psd*�`ے*����xB�W#�'n~7�bG� ��1�ǘ�1o<�4��ґ}�A�r�0~@�$4�X��|������%a�qW����&JʖRuv��V2cxs*�*ΠU�wr� b�*Rh9˓���(-�m��R�Y�̰deȜ��<��|r��C/F��E c�������9�,��H��y�zM�}f�FZ��W�q�d�7"�:E���A��'�C�yCKΜ�?]��P|�,c+:�o�̫P�lr�8�������|�v@7e�ly1��ǳ�M���L��v��J:�K:�6��}��r
�2&�W�堬Å�γ�AV2���<v㓷?bܹ9S���GR�x�$�F=gf�C2�y�]� KX��2JMg$0��Pe�dcN���z�'����kT�>Ō�(%��H��n>�����5��	�7ʈ�r�\fsl�yMZ�ۗ�*�H.D����x�����6 (cˏd�D��x�J%�S}��+�-Er@�ܳ�����m��Q$0�
+:Ȝ�b�G~!B �6�ʍ�8���1,y,��"�!��5���q�]�o��{���0�F3�ז:��N8�b��W#u�9�ш^-������JӐ�o�@�y<���������(O!uت��21����5Z����%����f�EIWdG��X1r䡕�MD�9�>�+���v��YB���ɴgP9M"���k-nrSu&���vR6�pV2-* I����r�WbZk��8��$�>I1؃Ȑ�HqG������l���p��9iqZ.�����+zc'�£xʊ]��Am�� M��֢�(aDT?Y�a�����Eȥ�;Oaj��f#lfU��b�&>C-M^F�B����/9P��E��0�pK��ʤ]�6����/1�~5@����x'	���#K.�ů0uWLAJ2"��X�q��� �T!9r�do�H+�J(�rUVf��ȁ�4��7*(ALd��2��P�e:~a�Ƥ��EF�Lx/�cV#�L`�%\�E8�FT����+�lflJ�2W8�dc���ñ?,`�V-6�EI�Z�/�y2��f���jB�;l�,e���NʥڨL��X��k&��Jpm�� �,@X�Pf�О���5r�ƹ��\��B�^��b�����(X��������ǹJ%~kfe.&Z��Rz�����&y�G��J�3O;��-WM�(���5=:Y��4�\���d��%|90ב��&o7]�c9޿g��9٨���N�SM.��{�*�lV�?LE���X��'ь�x��Y��گHj�K'̵K.����a�):��e��2	n*��(�X�1�d��(��������yp���t�W?�'A\L���0� p�ԁł￵{*O���[U�<r�����2:ta�e � <�-A5k0���T��ȋ$r#zd�7�#L��H���׳��󹝫�aڞ� ����i=q(��wNb�l�ե ����>>Lx���������*�ޑɧ�]ÿW��T�`Q��$�8���?�,V�G��;�g��!��^�QXǠ��^&$�4��4����S��=,-M3�o�ϹΔ�ޯ��.���8�n[��F\i�����VK�i�j4ƦD��	1�D�@��5Ϳ��]�f���6�d0�X�9����A�Y
ݲ���Py\֝�6��z�oI�4�;;zSYE,mV�+*�10$O!h��������Ο�s��y�tv��N��?Tuމ\+��T��t�S-5L|,�-o1�a�Mroƛ�cj�ew`ڼ��WS�iwe]��=y���29�o}�Î"]��]��ڭK���t�ѵ~Q��3�K��4U�� ��Y�3?~��)T����ˡ�7ݮ�����z��A�m[ꎡ�zsN�zxj��n.ma�t�Bi���#N�l��&|���N:5=g����ٵ�-wH�2x�;����4�S��3�����X+2,Q��܅�R�_�z;\i���i9��kGnkxaU�����y�c#�H�[��.��3�����k�4��-'��-#�:��6���V�=C3G�nT8e�cV�fL�U�|U��$�Dz�tؿ��rn��C������x�I<�Y�bP��$�"D"X��{;>� �B;��_:��t�Ͳ6��T�/=h�|��$^�@���I�I�Ks�z����K����9}u='�}�7�{��a�'O`h�dh�]U<�aU甐��;>�,e?U;%���:ۨV�5M����R�b�y,�rH�$A�(�-`��F�#�;�_F4Kh������$��0A]��Ld�>L�%�$�/�ƃ�\�����GPҽ��cV�='L|����ͅ�h=3Z!�>����t�8���9�̡dح?�f���,��z��+t�N�����z�d����;�Q$bG����v���u�Ř�I�{�%���U��BO[�#.��18�/%U����k�� H���9�?�]{�˷���2��6�M�K.��3?����=3)�.ZI��Tw2Nup���|L�Km%�J�-�����:��=�I�ʕ$v��~�I�-W�k�۵���]b�}J����Vn����*���c�p=� ��{����a�>�ѽ�t6�ݞ���+���g��m��u�m��wM��2u���I�� ��g5�?��²�%sظE����WXj���k�� پ��c��z�1Ӯ�Ѻ���$In�7(���C@�׾�[MGxUN��*�Ɣ��Eatf&#����̮�Q�c8.|�������3�7r;S�,p��5>��z�}��+�ҽ��m��.�t�u'�;=�m�t��+�Y��x��U�i�P�<�m��'Y�OE�Vw���gD֫ƞO���4d�B�jo?�������V�N�ݢ+�</�ovEQ�2Ga�\ӥ�j�7p�xOiU,�4���ctF/o�w���_Q��c�0���ȶ����r:~O��c�|��U.Q��rZ���R�%�:Z��FQ e�	fS� �O� 	�>w�����o����� �\ މ紁��}�]=��O�_t:C����{�ֻ��OQN��6�n�7J�楈��V�'S6V'�{���8�G��ai���L�Y9R|i�^Ы��>��k;�U�m��"W[q?��#3աeVC%��)��p�J���!���n�J��	��5(�@�a�Rr۬�`f$�Nb%T��T�C�'�~�v��:è� L.��׽�?Aga�}��v�;���1�NP�M+�Cu������M�:Ν�KXl��+N����9"HЪ��.����=������Z�F�O��͹�Ry-խ*��HI[�Q�NF:ֻ��6f�vv�P�S��⬶ >T���#A-��U�RL�4?.ǳ�vO���S�w[�B������ ]k�Α�λҫ���'R%���K�;�#�b����Գ���~b&�*%#� ytkN�p>�ѽ�5mF��K�|�z�Q����Qv� �ʑBN��!�A !���:���ҥҺ�����J4����^�$� Xe�$����Oi�=:i\*-w!����f}��6��Ӿ�� ��ݭ�����o�ܴ�;���� U똦$:�ܗP6.��wKT�ik�m��#Jc��X��`�w�d��ѫ�z�݅C��)�k[��l���G��J�P��&�J�,JVĜLxI��]Sp|��5k�RZ�T���]jXU��zi�}N�"C4q�uh��=����3�����+���&_m��b�I�y�cD�ҽ�{��\J~;w���9��/c;��yOW���蹯7}SNŶ,D�o�6��ؗG���Hj�8�N��b��i�}����oY�F5M6;��t�j��?��������N�]kZ����Wm~*F����E��k�$vd���V�Ӊ��V(g1{�ߑ�guV��v[�������;�����u.�u�7��{X���[�V6"`k��YieΡ�-�`Q@�����ܷ����g{��0���r�ҵ
��j�����G!�yk�;�6��E����j�L�9�障C嵍>���\@�Vz�GV� O�Ɠ������:o�s����l:s���{{��]����:s�ڞ���XZ橤�5�o_��#/&]C��%��Ó�Z���Ū���۬�#����sb��EӶ�����>��е�Y�����^H��K�e����� �T��'�,{�@���uMyD��֢�Ye�\xe�H��<�YJ����W��zWx�)�~ݱ=�v뮻��[�}����w�{���?v=���r�Lsp�o�5�C�ݿXj�^F_Nu�X�Pd���K#sH����C���lt�R��h���24O�ַSB�u��2��h��M�|bA_R��
�dx�I��O�����J�妗5�?k�u�n�/U�fh��&��p��c2�w�դX׵����x�Ӡ�G��e��}�������r���Pbw��X׺�jZor�_�u^Oi���3j����d���3G���&�k�w<[_��wOw\��V��N4�� 
M�^J��7��R	L���H�	6������۶/�mͧ�-�MTY�hO������M�<�*A�]%�4HҀ��6l�n����{��C�3�;sםu����F�J����V��4�W����r'k��et�����w��|����:.�gT�_¾��zq�w�u
�N{5�	�EĆ�;}ՠ��F�Z�d��y��Y���W�(|Ih4w����`�ZXf�IR����ye����K4eD\G
D������G�g��ѽ��W�}����.��-;�7p��ۯuz�T��`kF�������W;���m��hҳ0kygp�RE������w&�ovj���-,5�Qj�+j�Z��׳UN�D�~���0��8��n���:=���Jz^y$0G�M�z ��r��0�BB�ߠ�Y�E�d1������q�$z����OC�#���>��ÿ=�톣���p���5��w�������y�Ǘ�$�
�� /�r�g�m�|9�WdnD�֎�VJ�$Q_vi	2����ĺ�^�m�3q��>T�qą�P�޳o���W���]/Z@�m��59&�T#iz�B��Q��Dv{n"��]�_f�����/vߨ�N���x���F��t���� �S$j87�'M�]5��l�8�ꬰ¾	�Ӱ��ۍ?*�B��Uuj.�l�E�R��حEu����lZ�E�F!�嵐���*�V��:q� k�U�z�� ?�SQ]<G��‎:�S�*y$%��	Q`DJ���Wݷ�� ԏ�������r����M��E�i=yڝ/E���<.��_!gԙx�1�q9d��M� "���ᙱ>������ZZ��Jޤ�J�j�ۂd��a<2�p�?��7*sx���=�CE���ujt�%)6���{W��T<2� g#��uS0����+G�X��-�4�龛G�_��t�M���tց̾�OP� ����=��>���i�_��̌�b��%��:,����#$�� ��U{��ֆ��m$:py"Tw��A,��$H����j�Ǵs���u�Ot}�̆F��=��wh4}O�24-b�y}Sb̺N>5qBG!���bP�;Lf �<ޛy��率6[���44M��'�ʋ����`#�R#�p�������6���GL{p�״ $a-v3W,�2�d�t��=w�#���jR_~}q�'����Ǳ>��Cu�WC����2;-�Z@톀��`jڦgr�Y8�K�h�-��nI�a��yAv�\7����2쵸��kp�U��̯���=����т�7sp��gi�nmR��e���'2T���ʢF�O�ojw�� � ���X��Nv[�{���SL�����\-o�u[j��MisӟHǮ��N��#ye�����L���&=�^���.O����.�%�a�hb�)d�YHI����PG��n�`�$c��ҍB�z.���U���,������g2 �%R e�ت�4��~�{m��u}�~��.�����23����t9��~���� �v��4\�oVϫ�5�Yά�U�=��zk�n�;pս~��4t�Ȯ�H�-�o�C,P�0&5���D���]G�v��{KӮ��=˰Ȏ���QQ�b�TA�y�����k�������ݳл��ѩ�S����e���>7D�Yx�?J�]k֚�����m��K0��� �c�[OA���KQ�עӴɞ�U�Q��g�����ԑ`���� nf���Ɵ�P��t�.�P��.ؑ��H"�[ı�#a��~�<��s���Oo^�5��=C]w��&6P�1�֘�K�mwl�i�����	��⋆m(yd,,��f�f��:\�o�*�;�F@�=���2G���=�#��E�(,	k\�C4�~�Pr�����s��G'ߥ?|��s��������5>��zS۞��.��z:ê�Ӧ4�a�p�q�n�`/,]b�����n<�5�DV��H�����'�jpd^��O�jq�ZE����PC�2��FFzM��)�J�r#�{Aࣩo�q�hy���_x=ҙ��S���]-ڍ=�	j�G��7�_u��f�M'(�#���#�����C��5�M��eUJ-d��v��L�� �W�BD>�O72O*|⮨�T��>1����9�ې??J��z4�Ԑ ]�}@�Ul��x�@���.�����A���� �����R����%�U�w܅��������^A� _��Ҡ��9D���ܒۍ� �� ��CB>ߑ� �~}����S�� �Xo�;� �����=}���� _�g�'�8���~�i^FR�8�ES���[}~~v�|����<� ,��\`�dY�}���6a����T|!�q�� ��ӎ~���� �+���Y{��-���.���_�Ӻ��_V��mU21%lW�����],d����'����Y�g��?KuM�{�^��O����i�]юKE�B��zԄx������m�n=�KH��L���간�J ���}��8�r�_��C�I��;/���z�Aw#�?�z/I�.�u�L���}��>��t\�7O�x�e��U��m+�ߘr�Q��jҶ����(C�t�k.�A`��Y��oA!a���I���v��폔UX%��ɸz��4���I��IZ�+�#�	�[���*IH�ٻ�/������[���������_���o-�F�C��0:O���j9��SH��)z	7{J	�i2�����#,�j'#�j
�iH��y0D}B�����hr�Y��Y��픍8���\}�x�sfR�?{(�a��x���,:ҚV�����-W9瓓���+�̽F�NKx��5Y[�vm�z�f�kKb��b��^I$b��ǖgv%����O뙼0�^�׉`��G*�"(�Q@TE�T�3/Av�0��<�=ɶ=G��c5u_��b� O�j��¼�j芞���6/B�� ��C�>���b�c�g׋�4��||[�Z�[~D��}1�{������i����5���Fm景�bZS�T��\��;N��ގ�lV�������f-^o������,q�Q�a�^mPfd��(��rg���3�ڻb��������ϖx�Vt1!�_�2���C%��
2|r��l�Kt���C~.L�Tu�&��Ny#Oq���Vw����ٌ��D��o)�>@�r�^U*����=��������~$�fiӰqq���b1ޙrJ�q�}����)  ̀U�~<X�s�%1�q�*2���$��~����9�lv�9�!ϓzc/0e����RO	��Y'!���6I��r~ �8�]�ˡ\�W0�4����p�.�6�1� ��Ko��ܝ��Hѹ��^5)��X�5�¿�xј��n^jY�h�*�l�K}�T���C�ֵ���ǌy[p�1�&����ũ^q��"���j]>\����=��>}1��XJ��d�ʎ�I�l�2�q7t��a_� �BX��2Udj�BY@edF�m����V�x�1%	o b��ۍ�4ڢ|q�x��	�5�jU@���.X�B�,AeV\��0r�����h�b�Wu�||�=1����
˜�RS��gL~3]�^l���X�6<C\�w!D<8�(�6`�a������C�)Ē���1�j�u|y�ՖB�6=x6�; /81ृ �_��;�\g��z�d<K>H������@;� 2�f��n�q��++�4�*�3>k9?ڻ�U �H���JX�{�F��M��g�d��l���X���y1�o�@�PR��ۉ���>F� ����6;�~��c"5t��k���,Mƛ���c�O�m� �� ��c1�)�%&* [�wf�-*��"�C�I���~��Q��`�H���	o�X2/'܅U��%Nޘ�<�)�Ǎ�5��
����+q?'�ŉ�݌�Ǐ�r-�Fjyrl6 N ���?-F�����4Ȣ��d�퐡���q�4/II�&[Hr�e��C��p�rMcTr�r�lɌ����]��a��P��y��%�LB��f�Al|��<�U�C��~*
�bG�1��WZ�E�{�D�h��{��t,�(_��z33�"�|�����h�d]�Z]%I�T��c͔��_���d�����V�"��U��V�Ō��7PIf$q�`W�$Z�T��G&���hY3�U�^,�N�m&kD4�zc����)d(V�I���A�>�n���c�Y���2��N�L]�q_,��ڼ�Mܿ"�����6nn���&�B�r◃�>+<�J�R ܳ��Ic	A'�JX��\eJIcX�[S+�df��gMؿ �X�#
�ߔ�ka9�fb�U��ٙy�%vf��� O�cSƊ2hI����<�i�2S^*���1��1eΈG/���	�e��k�u�V4���I@vY�f{���ǑGZ=��¦���@˜�#�TV~��Lc�Ѓ(��	�k,s��V�)8�M�����j�~w,`���H+!��a+�[�dPgb�v�eJ��qe@[�B�1"<�Kդ�B��)�4�S�5�^'d5)����!��?��Jť(����U��褲#rv> y�T�ı�`��U/zAnd�l��4�%(]���� �~A@(7��n��y�ؙdFKt�rE�%㙜ꬴ,[q�<�ǈc�&��ϔ�EM��y��3VFu^&`�
>����*�q�2b�=�Ҕ4����bR�|�4ٛ�nl�i�,գc���|��F8i����!9*h�`�)f�X�/40�$�X񬑔���_"��2<T�� ���ܱ;#%Lsw����4��/ ��4F�շE���;�w`�(�ı�X�Ԑ�O 5�e���2���b
(	v n�$M&6�,�����\�PQ��b���`�*�� G���Ղ��o��)��|�w�( ��� q,aoj��G�~I#�,waS(�B2�1V$�?0U�E�QU������E��H�LJHY��P����	�,exEg5Id�i3��K�Ǜ�I4����y�N�0�U�8���1�
-��B�y.Ӫ� ��(��T}N��%��1�l`��H�j�-b�G���a���3l�*�4�.3I�>�eH/�*r�|��������c�	N��[�� ���Fo�<��l̒��H�m�wf1�V�s�B�.=&���'|��V,�c�IQ��j�NGf2C�E�~=�" eEM�M�� �^HT�TJK�Ɗ+?"�EMT�L�|Ě7 �Q��	}���M���6B(si>T_Ƞ�3\�fS ��Q��PFİZ�cX9QJ,������m�J�ېc2�wVj�x�LdY�E#ʱ��j�j�������D�%BW���'�o�Kc�X� �����ǜ�4��G��� >�ȋ��qZFhU�Xn��c���8��Y�I�,�A�Y��.����LA�Ťh����Tr�㕧9�iA� u�Q��@��k�Zvc/�_���1�U���@Y����_�1EߓLg2{��7M���BMr�0���]p�x��+)L)��� ֈ$,�x9+|f3�]��٪t�fV:�z���jc�l���%�fȷ�NE���Kt�5�c5:-12�_*T\U<Ğ�r�'�L��aE���,�fj����{c����Wj=/�`d��i��6���ڶ�~Q͋O�+���>wȴ-լm��ԧ*��uE�F��i�_��	#�A���V#�ģ�q�ô�M��,j4Z���Z7뿂��ֲ���� y�+L>���g��e�X·�9��=+�n��z��ǞĖ{bt�QYW�k/&�C(�w8UnGrPWH��ۺ�~�����f#�M�(eg��B����������f#�!���� �퉠�v���o��TӢ��Q�:����/-~Gt�VRW>������ޓ�!����oE������J�Ti�F��(�7]>��_�'bA����ޣ>�ݺ0�ZשfEQaK)��!�BXG����Τ�-�)����6�m˳u��d�^Be�ø1�$C���E܈��9�=����`�Wս���c{}֚�Q�����7�8G#�+s�/tVT(ɑ��KP���Ӎ�-MkB�cJV[�f� �0���;3���v+PXv�rU�z���#��z֩0�����Y�I% <�	��e�JM�*7�p0o��;���]��]w_�z��t��w]iٺNFt.�ms	z�#�t����S�,���عX�x�:X�Y&�h�>�����F�,:uM&��R��ʶ�H�Hj�9UdE_<�ȡ��{�3s�}RMW��(l�
��Ž^�I{P�x����|���;�i>V�����9U*�z�����I~�ݻ+ێ�t��ә�a����Fb~�I�ގ�����%M�����0���q�� w/#&ӦCȎt��;�Rܢ$����r���\��� YcF=��G�"(�����3�="�۩�=:���6�PԭV��#����A�	�L� �%���\�4�{=m�>��p��� w��-{��s�Ϲ���\buw\�ƶ�l�����k-?�=����ai�z�?;*p��pY�����i_�=[Q����O4d,ǹd
����Ӵ����2���z�-�R]MӫY���X��H�/9R{�ɑ�c� P@'�ϲ���K�~����׫{}����]7�u�Et�G�Ω�n�ղ��_�����k�g$�	�4�L�)f�V�֭� X4=NʳTj�Pc����D�T�2���(1�Oa��4ִ-2���kZ5��#y"WxVP$@Hd�$�r7?������C;k�� ��Cܬ�j�Y���I�0�����m����޹��~�ꞐԖ�T�=�㘧H��1�,�{u��-^�|:m{�I���&��jΊ�ۛN���<�y#X�!d�)��H�g7��b>�uOZ��_���z�лA=���C�ITY���=���&�X�S������w��ֽ��
7�/��ur`��=?Ҙ]a�z���Xh���M{8k]'�&�î^~��.��c���%S��O�ZgL7����4z�K\����'����v'���}>G"5��a��|p@�o�wV��ݹ���s����H��hB��"�W�&���v8�y%Ӽ�=<֡��Jp�y��jc���������m����t�Wu�u�^����Z�!�h#�=c��jX=4������Vzf%9�`Bv��vmxw�S-ЗRСg�i=��`�%
�G\2��ܑ��2�'�^5��EԷcɷ6�k1i�����5�OW�Җ�(/$���j��.Y�y�P�s�S����_^��\>��g��n�M;χ�Uj�\���:t%�E��Խ�~�w�M��ӣt�t�O�sW��\�$F�l����z��_V���csG/�W�T��ܵ�1��+LPh�4��mV�[��NPf̫�=$Է˱i���Z���nMnQ�H�B$�;D�WT@�҅`���ܲ��Lt������uG{�؏|��wQ���5��._Ot����-��[}-�Y����F�K7�sU�qʤ�̋d4��X4ψޏ��i��ҝw�.�z��<Z���#�	�4Z�T�-�����Q�����@�~�о�h�jͻ,/PN�$w꿆M7rS�9��64K�aZz���|zm���,�;#�^��ݤ�{��6�:ST���Odz�G�}��z��p�t�9����݂�llL<�j���2\W��(�}u��Kt��6�ޛ�4͑��.d�Kܰ;I,r��MR�	*j1ʈ8j��7o�TB[����[i;:N�ӵ��}*&Y�錕�i�rҴ:Ν=��)��Ȣh5��(S6��]!�}~�~��[۷l���z#�����ݷ�z�T�΢�}d5	cw��qO6'Vgg#d���ƙ�v����^������=?�_�z�j�[�V�*�P��4z�Q��cM�	��i nyEvEH^#��Hq���>+�CU����2S��F���^�Ԛ��]ּ�#J���<��Om^��GY���?�gC���]C+�~��g�ݱ|��u.�H)o�/�����Y��z�L��V��L\�={�Kk�'q��WiizN�Ә�ڶ��&=� ���-]+j�gl��=���D��/Zw�6��މjz�������Z��^�o��5��JR9���2EeXv��S3W|���ۣ�?o�U����;��'������os�#����m��b~:>�?6��\M_ŉ�����#U��������wH�v��-���]�r��dm=���i���"�˥�/i�<Vj%����[��������=?�+���r8c;{T��� �pkO���I��F!|�Չ;-~�x��=��x����F{;�ע�������7�u���.��zrx��P���:�6�M;���_/)q1�Lq��O>�E���������}ON�2d1�ٻ�X�vY',�C����>VJ�Og\��Y:���kt�T��[�4w�8v�+�?2����Ă�W�'�<��ٜ�;��ײN�C��#ާ�-��9�k�'�����4��L���̦Th]U��_M� 4@˿��p�0rg�����k��eVp�Jk���շ���{^Ҷܻrf R��]�X�T.�,#$�ߝ�!��0��mς�tZw��R��+�jVz�����"���I�Q09�������K��u,l=�����}���p;O�w��}��S]�\��?St���{{q��C7*����C�3)�uE��͵��c���+���Kv��i�U�-$ZY5�Qx�՗J�$`�R�^�}B_��g�U�	�:�{���m8��m[�O==q+I&���Z�:�D��y'�z�5flZ���?�GT�_�މ��� �_i}�v�9z^�����4��x:�^����o����$����V9�r?�7Y,�XY3z`�g�|/tgO����6����gS��F� �j�V7ibx���~��I*;#�3���j� �\�{hRt����
VӵJ3=��b�2;Vx\����R�����{���U��]����jꞫ�T�+��稻9��vw�;o�Ը�4,���:OT��W|\F˧᰽]<�9�SE���{�kL�>��uKZf��g�#�{���6d��-�J�bn T�#�=�e�?�}������4x��?���K�J���W+yE*��,��������m�ˤ�e�7���R�Lw��Nr5�'
=�l>��x��n�ae���LmZQ��jj�N�a��O%�^��S~����I�?u���䎔�y����w�	|
�N �lsm�{+]5/ �U�,�Q-�£�]E�;��b�ݱX-$N�� 2:�������l���N���WTfe�k���H�	�y�]3�u�U��=/�����hd��*�w�~�=$�4�Z]G�5���Q�	a������0"� ���(=ǸJ~s�z�=�(j�nY7�I�)-W���3�p$���+��)�����w�»m��W;�8���;ѡk�W���uL�/�]-��Zn�����Ĭ�=R� �4��Ɣ���D�f�4Y�?�j����4��[ԵY�EH#c�
��/d����4"N{���J:c���]�4��<�?9��F�;c�����۞ �<���ϸ���������U��G��Oo��}7ֱ�l\�#U����r�mo�:�MÖFf^66�"m�V����ǧ5q���������bu�F���F��4wx���,�ʠ�wwld�O�;���,����%�
y`W(L�pZ9Th]�@�1���P�Fix�=E�����E/�2ҝQN!�8��K�P2ɒSŒ2;Wv�W�m�����䊞�v��~$��·��N��#�#w� ��Vu��M��k�b��9�1xHX�َE��:#:I�0���X�@������e}1�ӵ��=��;��5��;E�R��oOv��pu=a:��:�O��d��1p�Sl�D�N=��Y����5��r.�Ҵ��jp�Z�lm-z�d�����e���J���y��+�l���� ����n�46f,9��uG�V�,��`9���w��3���-;�����U�K���ۮ��>��	k�Mꯠuw���s/��`S74��O�:§7r�
Xa����-2���Hd��)/�@�"��X� +�l�2�ee#��楤L��+�JGE�i�Eڿ�#�C
��]�G$�.�������]�\��ν�u�tseu�~���7Rw2��&���i8��5�s���vv�o�Ŏ&�̺~]�����t��f�,�^WT�R�vȌ��#$k��ܡm��'tv[�T�H�8+��7qF}/o.܂9�a{t�=�v�C�s�gP�5.��d:g��7'�}ƿQc�P隬4��2���.�/��mV�#`�rʴ1�LZ��b�5d��Ul�"��}�Q��I絁~���Yx���Ӣy���_���D�����<�>���bx`8-��粒��{��kn�����5*j:'C�X�'�䴼K�0�f}o[�QҚ�{dgכoT�	�7���Q��"y ��jF <��ʿeP9�h�$m��^@;yo|/�U~ȣ���	�y��dn,���a��a�T� $�v� ����9�� ����œ&�A��7B�����rF�lϯ���� ���Ǯ?�-�D�`�q�;�?��n}~����w����,O�l���<�H�;�� ���>���|�ǳ�'1]�"�j�s6����}��W�P?���ǯ���� ���>�9?�s�p�����$~܉�qBXqG�Ï�A'q�?��(�iѤ�f
���;1
��,�H
 %��Ϭ�gTF��" ,X�  rX�G d� |���c]��޻�.�M#�z���B�[u��}S��Ibdbj�������Q�4|K�Q�S�d�������>��ݽ�w��٥oP&���s�m
��x��J�q>�7�D�q�#
�}��j�cJ����~ߘ��{j�'��&�6I�G�r	9+��\�2�w�G����S�=F���^���:����t��M/7S�fn�����fdfGJF�2�t�ҵLlt]�*�=��k���5�oCk�c��S��b�DHY���Z�T+H���s�|z-��N܊Ĝ���:�;�E��;1�� %*�V'��Z��Hŀ���_�I�>�uN��N���;k��D�N���	��:#'�j]�� �����H���y=E��{Mj�д#%����-��}��y0�}v�F ��+z\�C�qA�ů��5�KB�XԠ�k+q�OvTk����F��/R�d*��}H�l�wH��o���*aH�lǋp(W}���<Ͱ龏|y�l4�q�$/B+���@�'.Q�e�]
Ѐ񢋠�Ռ�M�0����[Ŕnד�\/��������7?�〳�2v��1�c�zr9����L���������Fɶ^H�,)��^�9F7Y"�V38�F�qӛ*���[<r1������լ����V\�0�R�RҶ���A��F3cz/��GSL�+j?�t�SSm�o"U�6��h��M�K-9�8Ѥ���ޜ�_Ĕ�m��ץ��ƹ1���.�o'�<+Tt�E<&_;9��� ���{��B�Sb):`�2�� �yN�" �KL�T.C�q��:..C�:�L�iL� Ǧ�l�V��{��Ҡ�n��&�}1�/K���B�3�c�9ޒ\�rU(���QJ�Yi�
��R�g�Ĭ\�2��!,s�'�0�~�`۰ڴ�e$�K� X˗��GŻ�� %��6?	���%�!���d'�6c$bK�%Ju��7�F���4z�;�Ƀv?��N���Y��y�pW�mi�Z6��j9�v�8�kG��El���b�T	6���8s�9�nt������Z���e~ٮq�T+�#�C;�R��N�-q��=�]X��b�V������rg5
�?�������PeE�2P���C!�D�T� c���Q��ḌLr�|vc �3D?�l����	aM���2���� ,S�oLc��5�,�JiV�1�!G�*6 !P7ӈ �1Ԍ�2���Y�F�4�R��S!\�@X�Ðv�
�%�P? ��VoR��Ɠ�8��y�
ɱI����}1����,'Y�.\ϒ���y�&H��;����@@��P4�Kn�tƪ�l�jԘ�� ��vo�7,?�1UޭIS/"�<`f�2��� ۈ��h:��ोL1Fm�1��&b�4TF��8�P�V\p����Ъ�E��fef,�Æmd[��y@͈���(��	.����nc�"�=�"�*����rT K��ro����� ��zc1�UʑGz;dl������U�o��&jH�!>?�]�������7��EF��le����l�@��.U�,d��.�̞V�O�ĸ��˭o�5�x����J}1��4"�li�Ɏ��a����i�t<��C�jyrDcJYw`fCe��r��BY����;�B�9�����H�$�k�o2(�]M�B�"<�-�����A%�ZR�*��(e�́t��h��(F�q��� ��a��)E���
��D��~*]x�J�$FR���=1�R���rh�4�4PbI2��>NR�$2��!��=Pd㴼���`�D191I�6񝱘Q�KL��ϖ��(c��9<r�ӮK ~�ި��Aa1=��bv��1,ʡ�C�v/<kdI"j�j)�J�Em�Tח ��ጦ�tc7�P'�$�ш@�<.Ć�vU!Tm�����zY�4�+;d�(���I1����ā���錢d��3�ja�	/1)�G�,�>%T�?ف#���W9ӑ-h�Q^h3}VjZ�(j����X�.K$�W�&�٪�h�H�7fw���@@��"�� E�����iҘ��Y%�f�2nY�9��*Ѓ�#f1��5����D�L����х��$T(%T' �n8�cH9���Ѧ��%@n!f+�^㕨6����1�d_'�YY�Z�dYyk�Ȩ��UT���u\	M�1�E�Y	W��g)	�)4�d�E�lS�f �ȇ�a��LcYW��gL���Fk4�|�9կ��f�����J�@��1aJQ%��F|���]��Aa��-�c#|s�����4H)&�բ2����T�2�)U��y3�!�T��d;c�5l�Jp*�v�geP7M����$~b���iBr�2Δ�ݝ��* ��X�2��o)��tI��{ j|H�QЧ�[�;l���7��<qh����c�+<1���/" R�%�<�����k��]Dc���8��u3�˝��c)ކ��K�+Y]B��`ȥ�W%��lG�.��2A�'�ʋ��Ф��fcnR[y'�,T) sc���>U{�2Q�iW��J�R��Һ�n���lʄ�c���b�g��$�<���cҔ��L�C*�n5#�c�	ğM
�B\C���`��ϓ���|� ��$�R�3��5�Nh�J�:Ѹ�K�UY[ec��� ÓŌ7�D���y1����k���~@z��uދ�~lb3\#��A����L�Z�+?�F<j�+�r}1����FJ�9�f���38tRE�s��(�� ���5�Q^�oU$'�����j"k��}�Ê�-�,�fȚ�O�jv���H�+�?�
���S�!v��=<��'G/JJJ1�� I(J�H�ӘE;(�+�q�
�;f�+���k�q�|�$�2Ļ��V�y3��e�}�1��dLT�+�JA�4]��L��]�U_m؁27a��d<�7*�@��CP�ԏ��f�v
Y���U��1qPEjIdi�����Q� �6�a�O���Eb�KrX��r�y0m�Q-0���no�.O˘��(eWZkB��3.<d�4[���������`�j��rme�k����f�����6��J�S���[�C+*	E�R�Z�.�6��\B2�ޜ��s�-�����c^��XjZb��ӵi���,�D������ �]���>��u��E��E��Jd�#O|Ǫ
���ҧ�Z�(B���n۴�&�C����tɲei�����Ҙ5Ǵ��d�DΫ��4�HTb�����d����ȑ�E�x;��o�J9S[VkX�����}�(�}1������9)���h�p��BUJ�R,�*~��n�I���>�?<����ݝ.�q���w�6�.��7u;[�R�6����Z"l���=����Y�T�f.����u��t�����i�%k�2N�c�#�K�ެ�z�e���ň� ��i�%�W�w�o_o�Z�nR��:���f�"���ަ��� lװ>�������^v{�y�}�HW>�z���&]��{NL�9�y9ةe������Z�sE�kUwf��,�FC�A�;�e��y�� ��R0�y��-�7-=�F}sl��ۆ&/V�Lyq�&��C���>���	����I�u��F�N����2Z�f���~>&�՝G�q��ԙ�{�dYx�4]�b�C��R	a_�ke��{���omG~#�!R�9�Y�d�ߚ��V�O�G
����t��D�,ړj���2D
��r��Λ������G���ُq99�'�`䶩�����=;��O���5���r�lL�l�,�?L�G��I���h��=�z�]KJ�JZ��d�[I���b�Z�j3FlԐ�nʯ�,q��ȧ��}6��4k̲<6)�ʑZ���ǌ���:a�sx��hwFI#wC�3�� � ������?��+������.��}?�a ��%�t�*�J��dD<�M��]/�՘$�n�f��&�Σ��o�m>GN~�>i�~���4��´�V�,����s'�n����5ǯ���W�?l��+�#��_��������1������z��r�]['L��o�h�0hZC�dq'3X��)ᕛSH�7�:���4�_Ԫ�Vu� �mBhZ5�ך@��;�3)�3�t
��B�#���=?A��� a��^�J�{1i�d6nݕ��/j��Gd0ƪ�K䓎x�ރ�|�w�����u��_��z;���SӵMT��_��`5� ���+	���q� Rj	H��]ye��{��v�I:�V�Ы���j����'uã� ���6%�����D�� ,��C�a��t����A���]޺���Ԏ�Y++G�Xꎬ�Z�Z�B���q~E1���236��tǹ/����]C�t�N�lt�k�[�.l}�{`��JX����?�t XOE�!��ky(GR�zX�sO�z1�C�iԦ���	KCR���{�^Yɚ̧���a��e>�(¦a}���]Z�~�T�M8̖�ⶕ���Q*"�kG�B�R�mbĄ�a�fv6޲��m}�t���cS�ps��M�M�S�'P�CB�7u�̉��Ζ�V��Kv����8�� Skx�N��F,t���zy��B��꿊AU��6�2t�9ԓ�������G�%O�����%���v�曡U�B�%�&F��4~+�U���r�M����#��	�.M�MT�/a����{Y_t]U����ζ�L^��~�tv���2���=WH�G�����MOGm[E�r��F.\#0I<6M9���4��x�t]� ҭN#�t�PP��ؔB'�����3�q8qbH�W3@��й�Y��%|Ph����;�L74B�݊�F]�z�ұ�
4�JA���9�<��" ���?O��g��k�G���^�{˨t�U���Av�;�=,�W��ku>��c4�0f��O>BKtg�UB"�_I?���SիT�z.����a'y"f��,I<�K'�Q�D/��:��Z���n���Wn%�~�vJ�:M��8E�Z�QG�YeQ<������}��ob��Ck:�����vc����m_S�<���OS����u�'��ӷ:�_K�鼘j KS�Ϝj�H�Q��t���f�[�:�ܵ��[U Ӆ�d�^:�)ĵ����M�v?�=0��ܥ�^W4���ԛ��^�vV����U �bͯ�^��ԍ/���,+\. *^uV��a�}�W]�n�ꎋ�?i����trt��uFj{J�6~�<� �Yݺ�5y&Wb:�/V�፥�ѺoT\ӏ��K7�窝D��{6}��5]Ϧ�QZ����w>�B�����v�[��#�؇�B�*��xV����Gw,[�U:~��/���]ӣz�-��X3Q��+F��Y�FW�N���	�@5���}�v��u�W�OZt�`l^�.�d�L�_躗Xu<s2ۮ�kL\-$i��kF���S��|q�U6�­���~���z$R#�QW�e]�y�P�27th󡆯�^�hݧiw�~��(��'؟��u{+<R��$��������(�{�U�UU<q�}��.�W|���k����� R��i:�w���s�m��.��e�7Jvk����L���d�a��+�_�luʿ����7���Bm/S�SP��U�ٗ^(��[��%kRxfy�bZOhÂ��Tv�h�h��ZQkRK^av�4�TCj���|��`Xw���}�鎔:>�����'�{��y~�;a��_N���n�L�?^����.���n���iY�'P��Բ�/��S'Pڂ�R�� Q+���V�;A��D��è5��=�(z�H�Ɖw�TG4BJ���e#����Lu��hj;����[iG,լݭ}n*�	Y��r2cՠ09�ly%��,��u-�zt�n'�l�a=M�΃��k'�i�m���� �^z��uJ����t�~&���R��W|�3R�e��9�R��V�>\j|�]cyY�w7�Ο�4c� ��$�30�eH����{+mF �q�8@Q|�~17�����t-.��Qc������[�,z��-T��̖`���{�17�]�_�[{��cܝ��n:M�;F��.����aO7;M�o���9�.ygԾNf6��i�6ḛ�y�O����SۑG�n=U���j�q�kV�(X����V�8'ۼ�#����ͣ��^n%�{��O@�e����PplM)Qb�=����%�쇐"�e�����3�=?7�w�os]��.��pN�����s@�m6�z.V>V7p�=�1����6Y��&���ǹ[_Js��7��>�k-�H�t�"�T�ڒ��IRh呢ԫ�B���/�ѩ��(�l~��MN�k�m�EJ�mǩi�3r񹇰5;�x��B�@%��s����gb���gRwc��j��g��-׽8'܍zV^J�;��e^��Ŀ�)�;��+A�w��n��{pG��-,C��D�V{PCf&@щ^��ٔ��n	5��^їmޥ��O�N�5I�U�ܽ'1����\ƒ��� � If��s$h�7��t${[��OC�E���a�#K����@�� S	��/�t��6&��'?;2*�_ƿ�l�
�z�m�_A����q	�r�%�οG����û�d�y���=���K�ͨ�󉸝�2���^_���y`;}��V�+�� �a��K�_h2;��Q՚�{o��KķC�Ͳ�n���:��Mw�5;�1LL�CJ�h��Z���H7�����VmZ+s��[���e�R�^x�ۢ%%'��J�$d�>mmJ2�F�OF���	Z�A[�7��.��O?o#�yu�4���ngd������k�v�ӽ�Ӻ� ku���9e���մw����f���zdC�Hi�X�� \��oP�EwX�'z�*�&�W��u���I,��Vo�n1�6n[��)n�6U�!�[]�1e�#�Ղd��h�]�;r��"��kQ�:[�{��^ӵ����c6#U�;)���?Kt�Ծ��՚gNh�t0�WƆ-k�Luʴ�&����mmJ�Oj��[KH����7��W��4�"��W���<�"Y;���r׭n�;����W�]oXW�q,��0}O �Ex���A��[��}���{��y�N��F���-+S���/Q�5;��]cB�Q�F���U�4.��ҟ"]+�c��	2c!���:#� iu?�[�S�"��jz~�FF�l��3I2��!�h�ʯ1�o��3�Ͳ6n���Z}?U��ē�U�����$�+q;�B��o$c�s�}}�(�����tZ�D���i���};N��5)>NK�&F��pz�	�%��4�]��%��j2js��QMP����y��x/�R0ya���Ow�Ɔ��
�à�S���q�H�eU>_얗�Q������m�~�7d:C���wqt��O�߫�:�G�z�I��r+��#Hl�]�*X�+�]�r��H�6������c
wĮeYd?Qd�o|eX�&vOE�s��o_����0�nLK!��w��}�/2����A����t�o�;�N���3h��E�ؽK۾��l��ޅ����]e��l�%�O�R����(�q��dܙl_��lr p�~>jU������zy8=�Ҵ
�c�L������\�� 3�|�_��Wu����i��u>��j����uF����}cP��B�z�g�y�I,(~>#S��S�c3Gޖie���7{(��{
�8EU��W����"�x�bI��$�O�1�<��z��<�5b��5�4�m��$� �C��א^@��� �>�<q���㜶ے7 >ۯ/������F������ _�� \�$� p95+R��TP������n@ � ������� �? ��� �� ��U�J� �W�!�`������ �o_>�<��������{�� L.2!Jl�>.k��)������ �_i���?��� _��s�����z�#P��m'Q�����Z�Z>>.��`RS���f��%��2o�%��ɞ>4�wI��������4�B�&���r,Q�����X���i
��fo���ھ��Q��jvҝ:��Y�ݣ��Ԑ�H�e�9bO<���?� O��;}փ�]��S'�un�����k��\h]��ln�Ȧ���� Ft����[\��L�j��ʞ3#Ʊe�����:->��h��n~��ic�)�-f�?@&�[wG$N�4���܍6�׺�j}1�.��nx�y9]B~���*�رJ�V�'�Wꀳ(��^���{�GM��N�tMo�#�PtGd:[.X��:aDh��\c`T�3D��f��Fc��f���$]jx5+��|�m]�X�E��}��~�pµe࡝�����dN�Z��[g��G #��R�(9n��V�q��Ջ;7}�bC�|�����t��u�֝g��������ԭ1�O����L��zɞ���B�M��/wf`����:��$�/��D�kFH� �)$���i�-+���/ۛ[I��,��Լ5�~dp��HbT�>~��8� �;yl,lmGQ�!�X�R�D�f�*Q�M�����F����2z�3$���:u1se��C�&�fx�_�^M��W\s���p�����QG%���%���M*��1��2쯨��?�aT�=��~+���o@]��Jf��G��fN����c��N���7��Q�m[SJ��]k��xΖ㎓<�Í����9�g/Oӥ�Z~4���O�6���6F\)���� �d�����q"1�?�}+%�4ң�$��l����5�6�L`ԾBi�Yrdd���3c3WLtf�cP>o�	|�l�ZYOIb�ň�K,de✲�+K)F34h}5���q�V�<�K�22r�j�\cE�K�խC�o��qc2�Oh�����4�[51ђӘ�Ȓ�2@v��{�?�f��?�rJ�rǞ>:R��'�-���#M9���!_Lg��Ua�>p����QS�ғ�#������@č��e�[P�O ��c"�J+���̽j|����> �+錑R8�c��O%�
Ȳ�'�U��^to���Lpődc�m\yV�Gȼ�i-�zS��I%��Q�>O�0�;RsW�����j�*��ZS-U�u
��?�A�űjA�-�Za�L�>�)���h���� �Aʀ�'�rk��E��!7yҌ�;�Քnx1�� ;�v1�������ݑC�WeZ�R,^)�y���V��Xü�JYd�h��pGz��L!�e�Om�ex�܂[���l����)V��@T4� 0`7G`����c�+AY�S�r1�Y ���)T%"kUGV� *�a^ xj�"��tF�H���<�|k����qP�o$@��ͣ�ư2�|ukem�A��.�?�f0��w���F�Z��坷ޣ�ʒͦf<ySfb���Ջ9�l���9d�#��%?��ۋ�T�l6'�z�ү
̴h�ɟ�-�2� d*��Ḣ� 6�}~�NlO���f��$��E���v'�����ݦ۱���#�jQUWy�����:]-bY��Y��K�1��p��H � �0 ���.&�������yV����B�6���Y���L�W���b̼� �cp	c#�Q�{ƴXӂ��[�Q��5�`X��l=1��r�V��� w�~خL���M��rʀ c�n���	�J��9L���H��!�Մ���X�*���(�GB�iq�Vt�|UyL��|���EUBIcWj�`�U;�w�2�U1�� ��1h��G&i��T�%C��E#�w͢�吶1לWu r�X�ا�MC�]��F��D�a�����sڒ�-3�`h*���2��?�ʌ'�"?�j��6/p���uW��� OBU��Tx��>.$ϕ�b��l�ƃ�v��@#v1
�,�γ������cDB��ej?ځ�m��^	�|%7��2������� ��^����1��y3ך�wn*��`ZueU���Bҭ�	eo��f'䱅�L�2<�9ڿ��[���4�#�,�7�T�j)L`�ߌ�R�L�֓<E7aFU�=�P����bc�5p\J��Q��j��~�	+g�!F����9� ���Eb�&D��V�ml�nwaB8!�o�~Cc(y��:]�:E��\����,�L��۲.�05���j+%2# ��2Yl���gz��R_�b?�I>���[�-�R�<�Q�)S�&�����<>�� �1۬�f�w�ދ6�3�vd����"���ͳ�*7錡?ڔ��(�	�\ց�k�!�Ur��4UERy�1��!$HУ��$��|h0�~oس5����*�;Q�Mq'w�xϗ�㏐"N�꣑���Em�i��
ׂ�|!Fv��v��^4W��9 f%}1��\� ��W��6h�Co� (�s�\΁g��uK��'�XLx�~\���L�r��nl��/�W�⥌&3;מ8T|P�(0��e��y? �O�V�����������rkiKxvUŵy������7;�.��LaTI=��>���'�s�5wRm���T�9Λ��lp���@�XUi�д�N7��f�A�ۈc$����Qʟ/�tF��q���RA��ɨ�UPva��ldyΉ'\�=K�V��t`� )(�P�r�
+,�� ���~�ɨ�w)�jJ�op�#Y�b�t`8��I'e��"��$�kJ��e(h��:	ߒWdf]��� '�HX�E<��:c΋�)O*J���^e�J*��ĩU
ʹeqə��ꨶyH+�3y�q@�~
�cŘ졏�1�*�̼�#�C)
�Ey&��4��D@.�f�v1� ��m���t
���{3��^Oχ؅�9G6c &�b�ٱ�",�w�q)"v�9��Y�ud��<H��c	�5�a3UL�3q��v��+0V��]�a�؟�Lb7�n�GzA�� Q��K1jqV��l�5~,�X�D��S ���t*�1p��io6�[`U@�3 c�;d
�@�9�&@��l��U���q��O��c�����N��y*��38��p�:qVsˋ�H�V*��+�<)��B��s��7P��T��0FrlU��l\D�h*xH<��H?����n@;Pbv,c�p_4՞['����/����Ab���b>?l�W�*"#��\L�U��W0sZ�� Y��錃��'�<�VB��W�!�����R��7,F۷�0���[��&���@W�y�P��;�Hb/!��y�OI�ʅ1��6bW��d�i1��O��6�7$) 3u�k��z��	d.6Rc�p�ւ�³qJ��j���.��O"��sc���!�sj�I��Z6X�i�xY
�Vw%m4�����$�q)���q���Ե�#7.�0�<�����HS2�l���������^uU�E� ��h.��y:.�y�f��|(�B+p���Yl#�7�l	Ir���z����[��:��z�Q�]s�&N�_d�vlMO��R�l<�DdP�e�/�wr��OT�Zۚ��N��$Dp���T`c�&��R��� �ϼ��F��{�F���^�_^�n{;��ȇ��2}�h�%C�\gg=�~��+-w�{�ؽ�ٱq�_����3�L7O�4�05/�\(��������ԭ&=v,;StQ\��fB8R���d-�p����=���L�d�V�访>������l�|ƌ쏩ӈ7.i��*�؟M�� -�IV���V�5�iI�z�Ku�K6<��'Su�t��YѰ�p�9j���2��=a��CP�nn�V�eK�)���-K�9����X]O(Ð�4	v~��c�3V�WR�[�E�Π���h��#�},�!��/_I��h}��W�p���z{C���L6gIf�:�3cE)&|X�dP�g�o���m�=]u���iqG�W֧����AܝÐ��0��b��}$���� S���~mP� �7<JH��0I����ʢ�l}�
�'<:�=�s��]ѻe�lΞǟJ�X������ZnFT6d:oT�#`땵�W)l&��~J�;�z�h�M:戗e:�Sr���H�@؉_�Ո��wFÂ�kڮ���ڤ%pQ���N"�;�Ҵa%���㷇���|�v��3ܛw3�=��{I�Gg!��t��"ү\u�Tu^e0�K����G�ޡա����򦝧`g��_�Y�O����t���ͣ��^Z�lR*S�Y��m�|N�L�D��xk!�Wt�o��[�;���l�V5���fk2�S����Ҭ��pR�1Y��=��~���z�������Q����[�c�՝����-O��m��E�+�]��ާ��[+/[�>��Z��7��Γ��"�%��M�[�W���u?�2��]�z�SW�҅#h�(�����
u T��9]��/C�~���6��d쾚��4���+Ĺ4��YgQ�n�Y�]�3Z��[#����4��H�k�wj1��Ӻ'Si���M�]����D�o\k�A�h�ڭћI��͔�����W������^��-�&���U�I�VHa<��,�+J�~ݞI�*[�;���(l6��T�x�����d�Yc�a�{?uD^Oh�B�7���q{�����W;��������[�ull,�	��k����h�)���w���L�ӿ����͸5z]Nې��	$Q׸�� o��R�# |f�D�O��s��:i�V�5�Rl�ӂ�[���x'�$�Z���<G�"z9��߿k���K��u�=#/\��_I�#*){��Y�R͞f��i��ղ4����D R.)
�D>���~�펴lH�>ٱ$5$��ѷ	j����a�B�wr7�e)"r�sO��_��:���c�J�k\��|rb�h�����]	#�~�������]�o��}�^��݇й�}�랉���XĶ���~���
�f>����ؕZf�xg�O����#�:ϡn���1���mE�	�K/�Ķ$�)�Ddz��$�Y�Z�̨��o�u��㛥�t����n�EŅ����,S��<���L�M�-
�73�}�t�C{>�}��Y����꾰�S��q5΋���f�yY�Y�лy��;X=��Q`bM������W.�&��z8�v�ֵ?5;lK�e�D"Gi%�*��8
�f��$q �Eí�O��w�����5 ��C���X�[���%U-��	�n��3���׶�G�������?�:�������kaJI���Ҕj�qd�i�Y	ţ2\盃m�wQK��������~��-� �i�#Gx1'�|L��'��9�h{QЩ�Z���y�i�i�z���T�k5��X��G1�|����n�{����^޻��wk<�3_�׺c�t|�ln�t�����cy��@,q��v�����☹�'y6�y`�����Sl��`�#ڷ�W���q$�\�U�+��q�P��%{5_��������j�(R�uh|K��]�׌9�)�l�+Ol�A��:�������7��p�/ѝ���ѿ����H�����"�ѱ�C��?��v�����1�,Z�k���� �t�Z��Kz��M^�� ��I#��ĕ�Y%a
�s<�fV��q�������kU>F�	,Q�yen��R�L���D$NA� L���E�'��K'�ߨ�H�t��R3л	ߔ���뾞̀��~�����O�u�7ɮ~<2�<��\���;���ln�K��IٚN��G�[CP��:���s��-��B���byS�%{Tk��Q�4sPݽ<�z��S�Sz�z �>��݊�r�J��wĮ{%���^���پ��p}�k���W헸i�R�gi�W]����Zj����R���y4�\�.�������ZVYW�Ը"���7�ޟ��u�3�R�'3�3Y��ZZ���"�U���Ec2��� �[�|�߭[B�nX{k�!�bׄCd���H�K4<,��L��?�JF
����� ����s{'�>���k����5.��Zgk��|\���%�t�6>)]���!Y�hvY3�#m�НjX�~�㵬"F"��4.H��J�ꡕ��/(v��RNH{Ϭ��s�m;P�ঽ�����*AVwif~�@=���?E��s���vK�{m�[�7�=c���u2���K�z���u*Y��C\��~�2t�s�acX*j�uEB`���Oc�6��4i�z�x��A{%
b^#�i"��<��+{R����E���Z�}��kV�t��'�8�<����bYܒ Q�( ��A�N��^i��;َ���^ !@޿a�"]	ԝ��m7+"�|\�h�����B�	����~4�5l_�Qw�N#�V=^��th��*�w�;-,��	k�D+2ԚEi*M��V~�_�������q��Ch�cX�-=J�Ə+"����1�K���u�T�cr��u�o��}�ӻ�{>�6��X���7�K^�z::���:��Lt�禑��3��&@cb��IǐG�A�y_U�՞5�Y���hkȧ�:�3�1xS׍�,�:Ǿ��ލ�a�P�?L�ҡ���R�H��9��=�n����v�����^����Ei��M�]mܞ�u�T�,V�4�5����!��c�F�V0���]޶�\��n��[FE��"�2�/ƕ��c��:,�ݪ��N����v�ۏ��3U�^Zk�,�<�	�;ؙ���Wo��31�>���c���K� 鶋О�p:�5���W�5N�jZfoVv��r�7����tmS#R�������kɱ,���$yS�t��V�%}N�&�.�-�"�Ԛ��kj ~Z���dFq/���L{_C�"]>���[O���3ւQ�Yk�@�g��4q��_���{��ޭ҃S���i�]֝M�����_�����iz�wYu��n��TF���fd�:����/��v�MiҴ�,����0n�Y��߼gc�O*Y�hz;�Ϋ�B�
��,�|dR���R�ʂU�@_����9��h?�ݎ��V������L�:�C��<}GC�-s6Rk�&��兕��;�?!���
�Jd��z���WX"�☪v�yW�?$?(�p�e��_pC�����<�fG��+FA3(�/h�&P�Ib����t�5�ݷ��g���z[��~GA��?H�m�;��|,+�ˏ�j�
m�tI��BK�ߟkъ&9J����Iu�5�����
�>뽀����r�$��GfF�IX{��[�LA�_�#��A��d����fS�^K��7A	��v�������� ��s��=��ߗ\�1朂Nl��6����;�_c���ׯo�9� ��9����Z��܈R
�&v��h9?�v�����|�����~Z����~9(�����F�������� _��Y���?�����J���e�f
N�m�m�<�#�돿���=޽�����,��n����6ȼ��|�'�g'���$Uț��+��}�~�}Ď-�o�|�y}�=~��U���y�8�{� ��3&h=��.��4���-Yƽ:&�u�21�Eq�,�D�1%(�PL&�i��(��mҍ[��m�K1�SG~/ꓐ!��Ч��P�#ZR��h�yo�7f�_�V��XP`�-4��݊f�-'�p��j>�=���V��[����bt�Eн}�m�]'�t�W\��L� ��-L�`>1����ı���[wK��K}6��f��Z��Ւ���jQ��EP�K0�(ɏ�JI0?Dp�*����tZ���
8j�B+��Q��Gu�㕙L��$��*�����]1����t.Vw#���t�n���2�u��օ�:�&�K鮉ӱ1�\�o��5z�ӱ��䳆��w�>��4�t�j������^�7?�Ԃ�9e��l����*���Sx��jv��m��~]�g�����
Ԫ�����0�JD���(��r:�P׺�U�z����Q�[]�r�5SW�5���sr��X������**�U�߿wS�=�B�ܹe��G<�� �쨠*T K�h��*W���Jt��lqF;QG��$�fbYۖvf$��tNc����w�ʃK�9����hO�&��Q�2QO�nZ�*�&�ޓ�0�_�X�V�&L��v���!�^#�M��=&�)e��e���m*YQ�0+!��wǮVK~I��#��5t�Z%9W�9�ȑf38��O@,�)i�\���qMe��c��)h��>��(ʞi�Z�Q��_J����������5�����K�O!u��%�N������c�HҮ�X͈�.��;x����I�(�\t�;Ta�*�1t�� <���~fd���JZ9����Ƣn�tI�c�@YcJx���W�ϐ��Uf�pfv�4�S->ڎT�!cWE�Sɨ�'�X��l��U��xc2v���fj�'31���M�a��0��eJ�(r�%����4�d4�!����%�\^X����mD�o����r<��v�A_Lg���ga�K�P�?��p�>,L��N��ř�G?��*��y^���.$������J�pi�<�����T�1!T��r�c.�s�t��i��Yo1�q���'AJ?o� =Am��Қ���nS���Uj�4M��*?�@c��+�E.q���v�INU���Hry�� �d?e�c%�#����o�|)ԏ'˚�Q򻢖%��g��
�XY����Z�UQ�p���*XIn�lU��`�,`�5&����=�;:��t������r�pk� 6UNO��U�s3�DDb�R���*��n��S����L`�R�>3³�E��d�o���0o�ۈ��&S*�z�t��Qv��uj1I�2�b �9�x#�~Cp���ߑ�=gc@�ҫ8��<�F���UC��c��}B�1�\�ڻ\�b��{%Q��Q�5NL��x�^9�!�`B����bǚ�CI�W���6��)�<#d�(}�m×�1�W�Q���P�:�栆%\�u�(p
��c��rR�k�ewaw�6�)1EVS�$����ߋ�q��k滅�x%"V�x�d���w�Ձ�K�������"�x�Q�+�j�$B���� ��X�f�	X���J0��Z�VkD �'^`��w �c�w�8�`��~ �9�����H�'�zc1���.ZA-`��R�?�x�ۭHe$�IT$8S�c+I�:�.��������_��\у���ۃzc$��Z�o/7V�q�!N,��7�=y+�bJ �ʒ5"NuG}� ~qҢ�Glq�O��\���AcN*�Q6�b��9�O"�姂���UU�*ޘ�[P�Gq5�>'��mWGs{2�Rs� x��vv1�	���F8�	�@�S&���!���|�0>T1���A��|�L�#L���v�]���wTn@��6H@�f�#���&^J��[Ċ���r�s�����e%vV	5��dI'��	I�5��G&%������R2E�ψJ#��"��D���
��f�}f=1�,�����/�|�j3q��p�w��*�S0���!O�2�%F`�k���2�:!�j�`�����~M�r� c|aR�#F3�A�i\#�yS񜗄Z����> �+̀�U�g�1���::�,�1�:�'���Ǉر�Iy��;=�}1h�UZ�MU<����l����,c+:�Jp�C��A^��XK,����3%���?���i�Ĥf��cG(��\��7_�O�'��q'oLeqC��0F��(+�0��؅�V�˷-��	�P��WE�O<���]�������c
��J��wbg� ����1�*г�̹�q��&9h��q7	f�k�g�m�^1=�@(�C��^T4@�7��<�_�t�y�c�ng�	�\ ������T oLcgZ�"�:�ŻUϝ�B��?v��< Vc�����D�ԶC���VB(S��bD����T��A�cIѼia4Ie�Z4�eRD�'-ڠ}�P������عh��\g�0i�Ѓb��q6bK�9�~l	`�˶Ǉ�i��%
7��VX�ܫqE�U�*���Lc�ְF*�+B�R&�BV��Aȣ�3��RH؃錩�P���73J�2&NO"�I�eO������1�l�zҁ��MMX�;5k_
BΫǒ�;$o�n�)�Iǳ4� l{Q��GFڲ�/!4Nd)j_s��,Ō��k�� �݃��Ky��g&to���#q�]�r}1�[%耺͟��9�j �9՘Uf�4f����'�w�ر�:Ս��	"H6�tY��?��a���1�z	�h��v�j��X�Lre�m�s��r�B�{��d�@Ԍ��`#ɕ�W~ �vr� ���f1��_�ɄލTG`�6�W��(n<&�����n�T	��\9�4ݒ��5���S���O�RC�%yOg�5M+� æC���Lz&��	R��>�Lda_-�$�()7�)�Z��	+V5�I�Ԗ%G�ً1����I���I��3g�h�cŝ
(a��+0x��_�����1��W�B;�l����T @���C�����I�*��k4B�K�+v+�%��<�o͌t�YJ걌�IC	ƮY�>
8چ	�M��>�)c�nX�.�e�85���"�I1x�fǁvf}�e��;�H2^c�_w�Ǫ�	#,�>�m��@S07eRK��RA��`� DY]ãH�jr"�.WdA�,�4���j>:c�s�ݹ���*>���B��(9�1��\�i��J������v.?�5)���� ��3ҨH�TV��Yڥ��nmp|�!��P����Pv�=�IBߏ:E\���uFn!��$�l�s�.�$/��|�A+QNnnP�Z؍²��a��3�j����H2YݲƑ5t��Q��?
��2K;+<�r<X�B�b4�����<hʫ���l���ҴC�G�ǔljvUy�%���g){��)�S�&��r2�����|�,K*����H%h�.�_��檤1���׷�S�K�cb�����9��#��3�MrY���d%e�oB�jVwO��ߍ�A=�s���K��So�p@�p��ι~����oC�:WE�}O;@���Ƨ��M/�&��j���g(���\ɻ?�:�؎��~ܻj$R�yhyJ�%S���؏�OvD�駱&�Ư�\�g�	�Q <ݧ�]B�)��!K(��� s�8�g֘��Y虺�����:���yeiWÿ�­���L���۔���[��x:Q���� eh��;�I�\�8�a�$G�x��=�c=ߖ��`�F�߬;ƹ�鶫����ִ�g��N	�3�ϦL[������Vy:Eٯ�;T����_R�R��r�u�J�.��i��Nq4�G�1e��<kU,Z�-�Ƨ�7��ѽ>Q-ݢ���3��kXO%YcH��������h�a�8���t����Mm�M*q_Q� ��ix)Ӫx�䈷ݤYx
Z9��W5��̟���::6fo}�h�_�9c�+��=�n���X媐i�9�Qb`�(�NF�Vo6n-)U�]~"v���COpl���'�K�5$�~����-S�'!�p�Cb�KIo|8��t���륩]�f���zT������ 4jH�%�$)>�;��aw���zk^�4�c��T������'����솁���f:V�����i�*�jM1Ɗ�x]�Z^���h�������'����&�+�#S#�h�{;�Rk/�8u�K��y#�G�^��{�Bۚ�ߒ��td��Ħ:�բbH��p���6^� 2��^�����K�?�;���t;��v�LίZ��{K���ɗ�L>�v�R����b��t�wRjsr�M21�IT�h=?ܶ�M.�~���\)�F���+���lOC�����e�'����o�O�z�4���N��g�'RO��rL�|~�t���D��a_�?�������}�u��]O�9ٝ���T�]����7;�p�X̧O�M���¾��h��jɄ�~�͓x����>�vս#vUo�,������F��2Y����23��ߵcvnx���M������@g<4��]�n�R@�&�[��Q9.����G���#�N�dv�Mв3�w��G������Z4�G+T�4<l����Eh�c���RAb����s�tޛi�w��W^�M�EM//^'�i��P�CG?�1�ns��˦�� R�eE��jZ�4�bf����Xܹ/�v����w����q�ߎ��څ�w��KN��M+V�u�/K�~6J����bͿ�Vu�KJd[.1Dv�Z(��}U��E�iu��7@�bd2G`m#2�ib,��A�3��f^�kgG��=3Y��P��Ң,"�{�%nS��RB<���� EGOx��f{��v0i�k�:7��9�x3�==��:7^u
g�Os��M[K���ŕy��4��;҈�*���|O�Ϡ3l9/���h��i�Yi�� ��Gf��h������;I�~��eM�i�ƀ��R�x�;�Xr�僪��}-''�Fa�о��#����;Ѧ{�\>�Ի����N���պ�w3+�r��L�q1u)By���M�,�� z`���z���~���������S�x�%ż@�����-Jܐݷ�Y� �*��o��ǗnAO��a��~]����'/ �"�;�L*�K/w�{?��Sw�Z��۝3]���m3O�)��~��)`>`����Y�፧5S��<P�yR;�J4=:���į##)��rF����
��+0ÁΩο�����W�!����8n��'��̜rˍ�]��Ҵ���_D�u�J�>6�>���:Y��:v��6b����;3"��9���!Zx�4���j�ն��j�-+��ah����y��<�}  X��v�Y�Ĭ�ܴ���1+j�\�VO"ن�w,6�w�;}4��r��`@����]��O�W��}{����.I7Yi��X}�е\n��p��v�P_:.>V�����m�:xC�q�#MJ�Z������+pF�X���n�w���1	 -�_ơ;���x����b����������;�"[����b��
�I!����)���h�C�#��On{M�_e�Eَ��'SSJ�'L_��P���u�P��a��Ru�!\~����y���Fi4q���WK���ʚl��0W�^y�!�X8X�>�,��r�"���;�A��j��Q�5",4����9˲v��<���{���X=U����W��=�뮝���)����>���.�����jz6�4���K�� L��o�3uBd�~�75ilh� �l�O4,v*̩�=A�rɚ&Y}���ٱ� Qum;L��$�{M��H嶓Dѳ��K�x����ᐅ ��Fy_u>�;�+��1�^ᴎ��r�W��tޝ܎�j�1��.6�����h�m�yҼ��g�t�\e`V�铅xJ�=�~��]@Դ�Q�˶�H{ޤ�:I^heu����"�)��^QdX�����ibu?Z�Pj4��T�1�Y�eȯ��0�H�F1���a�1N;x�>�=��w�k�}�{g�>����]_�����Z�5���rƞ�=WPǞ>6��b��!b�(�`7�5kf�?��.�R�jMFKn�I��K4��"ݑ�q�
{4@K0�vn[1���-�n�Mp��h�"� �B����� �wrH(��������n��}��� s�~��p��.�T��7V|lC}G�u���\[kT��o��!��n���ж���Z�iD�5=D�$6�]�H�d�d�[��*����m���Z]]nВ���:��bU�3?<)�G-<lpH�ҞH����~��g��۠4���l���p�b�wMSC�q�&���/V���qc\�\�6�\�Q��ӆ?��%�Cz�k���S]�Q��,�*��݃�I�����>���?��$i:KOK�Y; ,���a�.X׍��A���|��_�ޠ^�龣�λ�ZN��-Jo��鍧��������1��o����6J]edCZl�5�5}&ɖm�q$P̝���x<r?�DG�	*��E�r��@И	��߹�{�%$��c�B� ��7�n�7�=B�5ٽ3Z׵�O�:���o?�����w|�1��G�6����U5V�sv�Q��=KG�/L�D���G#(I�px)ZTp�'��G��X��:u
��ʫh�d����9Y� ��<1(!\w�|�z;�ֽ��ҧ�K�:C��N�н�����}�Z8���4m�9����o&nc����{r�µ������K1ڑ��#��#�{
g�h;�F2M!�������} }*�>�����Mull���|{9c���7��� ?������?��y0!���?��,�<�7�L��l�~$�m��o����?q���g�#�����vf�@~A+3}�}�]� )� ��� �������� ?��?���W�%U�4 ���\�"����n@|��}����8�،��[�bv�S�ȫ�ۗ���o�~~}~��׿���~�~��2f2�E�U*�15u&�8+�e� ��B�>Đ ;�������� _����g�ׯ|� ����o��f�����5�����o��pza�a���[�t��g�i��x}C�8�<�}M?Dc�Ll��pd|?������s|�+LJ�6̎e��٫�M��	#��,�M/jII��f�H&%�z�V��Ojy/n9c�+1�IJ�ܞ��'-��ξ5Wb}ϳ���'���Vj���а�O��e��.j���[IҴc���E���uLM?l�Eu�e�|���-S~ꦂ�m���� {çV�R �l�ś2s�H�1�5�y�t홣Es�.��:�p&*d�fy~����!� 9,���4���������r�����~�u&V�ڽOE·Pk�U��z���s�wԴ�K(,�����
B ��2��a�3�֪�b��&���{��<�T�+ �a�XqbPHs�"�2���w�6ӵ���	+Uu$��ǫ����ֈ�ѣ��3�ݱ�=_QȘ�k�oŚ�!��g�mVI� ��6ug#a�~b�8�=����ھ��H�> ���1r��*s�-c፧:��^�U��"W��Q��.���'K�EL���C@�U�F�K��G#2����z�;��iyĕ|� c2���ej����΢V�X����:_76���N}G���̆��Z76�Ŏ�̽�=�̾.E'�GW�Te��1x���q}Bx����|�Ϗ?�u��C�$�͚�>��^6w�Ih2j�����~<-?���r&)�g8c�kȡ�sʋ�����;��DֹI�����ͺ�&6&V>@w8�ωI~S�y�h�y��*�7c6J�?e�ӕ��1em�^OVj:�b�(�mĠ�>J�;zc2���L$��b2dX�*.��;�Z�i�TC2�~F��L�����J���^q�'�_!Yq��[�c��b��pU⻕	���k��5��Kl��x��^�ч�%"�� Ls`��nl̞�����%��ɬNsu6�p�B_I�+|*X0$�۱��`�D�ί	�B�YP� ~8ƣ���gڟp�P�JF��t�Q�ݶ�xZ; Ei�p�F.v!��p4 �^p�4G����#1��f`J� r�(ر��Pg9�ƛ�!��x>BU/{}|tR�9.����by��*�q�+N,Y~�&�:���AZn@l v1�x�xxéȚ�f/z+'�����p	Y����s�h��:WX��eI9͕e��#�lW��c�|L�fUd��7��P��<��  @��L���}1�K��f���Td���4����Tf<B�@1�6�����1�L�ը�ƥ�(��{l�6�%���Z�FUV�*��	Y�X}_�-)m�}�1�-G����GH��-��U��~_�l�&���D�Q���#*����YZ�fe��V�pq�,>>W�pX�lvE�����VV�ph���ߍ��X}� $��V����|Y�jx�W��]V�Pf�J�R%�²�L`�W��q`�@m�������~8ER���W�cW�V_�y<T��75����n�h9p�1��r���b�LdP�j����Y-TQO>{��'�y�.�wřIx�W�hTynԖ���c��� ~���F)$�x�$�¸�0?!����� ?>��w����7�ﴯ�|_��y2�<��UCpP�hO���d�W�P2U��g��w�B}�C7����c�}X�TS#�?�s�c�|Q* *��R�D�ż�]���\)Fg�K�tc��O��	�
͚��?��b�}1�eU���x�Ix(��@�����%v�cȞD��1B��UtLb�q`6p(�)}��U� �rf��VD���_Ȭ,���HY�r�kF\]��$Ob�7>[�d�v�r��!v[�kjX�Y�[茎|�CZl��0n>/��"�P��!c�,V�"�Fb��6
�ClA�ɀ�CSC)�ە&�b�O"��7�3̐���-��VJ�뎭GE����Ҏ�+�*N�el����<�c�<��mـ�56��%�f�ѓ�*�QN�b�.��0Z�4O�r�?���M�?�$�7-�۱��B�����Rrz�A^7�gb��s�9N�W�I�[��7�r���!��N�Z-Tn�QP�� �c$L����t�tf�� 6,�Y�:̈r ���0n9���!iߝ�d�(	+_�9�I�Ǐ�O�,c$����E�7���F�Y@\�-`J������ ��� �B4y�J��h�̴�n<�蜝Wd�����U�lů,zM�H�I�wV�g5.�|1�� ���<U�x�)�:�@��|Lpe#��,`dM��Խ�JVRƆoe!b%�c��*���$��bg�"��B�V`����ڄ�~�bJ� ������ϓu�vp�ч)𡐝����n�J�~c�I9�:�Q�Ѧ� �r�ٶ��(������,b
��y�sh��Y�j�RH~ IX���|�G�7oLa�Ѥ<��-�HR4zP��Y@�*����@cf��!�LG� �N��Ƞ�f��qQ��G |�db��n,�xVxյh�\��BW`�HbvD�1�D�8�iӂsh�*�j�ǀ�q���C��˻s�1���M��n���>[���&J��
�,Ԏ��ǴR/@e���m9�UV��[w��f��}Ϧ1�uZ��M��eGC"�w��'#�,J�`C/"7<�āEX���9�ˈ*��UI�c�Q����-�7R�K����+�0�]&1l����Y8?�8��UJ�)P�`(��wO�V�W#��|R|�x�r%�������bK1|,��Ό��^B��q�eJ_�X��#ʛ1�%�M�+
�A��*���Ρ�oB@ �RD�`���;���_��us���D�����f9�į�I��c�����q$�v�e��TT��pImڤ}T1��TzKud-�^�;Z�&�4e�o�x�,۩ �Ǧ0a����v�yʷ�F����I*�U���x3�1Аʋ�/��KY֣��dK���F�[���dP��ۣ�9��IzsMUg&tq>doNy��[e��I�D����F�=�S��P��q��~���n�GٌJ��CH}���@��o�'7L6�b����ɹ�L�/-��x=h��l��a�(��?����B�R̶Y͕�i-�@O�<)�U�M�"���1�W����l���C,�q*,��ٙ�2�ٕ�*X� &r���<�"�|�4���m�3|'���2��#�4�q�ְ�C�Ƹ⃝��6�Y#�c�f��a�I�N[�B�0�))���P�Ǒ��f�zc�ɋm�ލsg4����v� ��]�k�n��;+'O/*���by�^��:���r�K9���#1r�fJ���f���
���sNn��/�<�4�3Lu<�c�'��-�1�c��g�Z�KMT6����&Uq�7,���x�����g<{��gK�'���ʂcd_$KL98�H��\k&IoSF�!i���Lg!���/Z�5;_7�����s�_*T���Uoye$��K'$���c�'3���".g��yu�/C���N*�DB����KO�A�u_#���˦�X��XlsV�MHo�u|�U�D�&限�YeզfFQ�:����,Sי��GFdta�2:�����~�<lW��յY�e9#�H䍇�F�Da��V�Ⱥ'���d�#�}[����HE���N�gi�qRκ�k^_,ةIĨ+��7C�/]+hJv���WU�v��c^���v�R����b�nu��R��%���e�L���O�L�`�B���e��Y'����'��hW�������hZ�Mc��:#�zo'��tZY�7Ԛ>�f�&Z^X��������ɒO&Se��~��W�w~�%]n�kܯ8+2w�{����>�1�k�1��0dfC����)��N7d:���&�Z�Up�\�4v+M��i�Nǅ�VH۽Q�������� O0����ۖ^Mu\���"�'Q�Zޜ��4�i\��rݼ�x3��j�o���P�n�Һ�Zƶ�o�?Sk�"[Q��Re���G�X�)a��b�I�
�]���U����+�<�ӐH�^F��D���q�{	*J��< R/�O�� �{��N�����z�^�Q�=SZ�o�U�_S�U�V���#�w��U�4��&���'ֺ^��;:m��ۦ�4�~{!���Jy<�iҲj'>�,@)'��Lz_��Ԇ�0��wW�ª��&��*7�9���oz�:=�O׺�����?����wlN�螏�t΢ä�X�ɟJt��\zO�k��ɒ��䳲���� Z��դ�R�2�^xO����!������rUes/�Pgվ/����"�qjV��En*�cPN�Ӌ������k0 g��Ow���z>P����R�P�2v�+�����:�RZZ���bk_��AA��ɼ�r���A�-B�V-��k�ھ�EU�h�I��>�P���$��H�� y�yʝ{R�LT�Զ�ɛR��HY��̏��`�jȨD�EI.C��^��A���c�}�u�oe:�Bc�w��I���G_[V��gh���jL��\^�vYddK>y�+G�Hz����5���t���4���j�E��Sё^�H��-����\�ʓ*6��b���(��ܩ_�sFlERc�n!X�����f!7Ҥ���O���ٟn�kО�{���ޯ����>��:����R��d�W�k}Y�5���^:���j �r�	u����]�܆����H�KB�`Geмld$�~I�n�ډ�՝cb^<횫m��R?3�95�0���C�whӂ��,����zy�n�ʿd�������}a��M�x2ƺ5���Ӛ��Mx��4b)J�Rf�}Sj�ԣMө�H��CM�#��f0�P�XL���*����WE���[n�^BE�/	JĎ�YfF�GF��j���]����?n=KՑ���>���ё��)��U�nx�C���jy���:/M�d�q�o<|�|q�"ˑ|Bl�cv�2/M5�"[��旵�(�s-yf��A�?��Q�da�,]����	���3�����s2@YP��v���k�B�R$��  ����?�'�n������n�{�辻�G�5��;;�ޡ�N���-K7/�u���ִ�LlO�c��G��f4w���!�Rt{�ˮ�CN��W[SZG���)W�"�Fv�g�(n։G�6uO�si�C�V�IRE�40�,Q�bc��4���X�K�e$���r5La��t������f���]P����1zk;?S�:=�R�y��pe\��힯sEV_����C�b	����v#�����P�I��R�o�$�2%��+/c�3j������dM���k�z�7K�1zk��G;�2�f�\>�i/W�mCS�n���_����������.CC ���ø��;��Pݬ��s�bHdO%9яtV;d��{yN�M�Mi�]N�Ս�FX%�ȍ$-�9Ae`8z��Kؽ�\{A�>v���zC�1�u֚�I����.�ѻ[���5����� ����X3�x��S���#8� 3���l����k�lϫձCL�f��x�K�W�rN�bJ貎����X��ӱ{��Iִ{�Ίj߿�J��Yj��3Eˬĩ$ƒ?��o,�x=��Η��cT���]W����uF���i�GM��>��,}R�J����S�9����y��Y����[M��5j������qr���ѳG�
żRy��y9�Si��[|�O1�U�.�N��0�f'�Hde�Oی���/����>��k�V�)fC#P�.��Sv?����T��]�Қ��"�=[M4Ɓ��l�	Y[W�{L��i��j~7�,F��e2���r�#��ְ�I�'�\Ѧ�v-F�h.������)�t�@=���<�3!�0?2�����vs�:��A�y�#�=}�}Z����}c���=s��k�M�=1�������9Hf�_���e��0V���/w�ܺ.�棪�*�ZhȵYݥ����Jc����ې� V�5.�ɻv��b�4�Ex���K�"0�E�9x�[�$^'�UfBY����{}A��G�����w/��*1�Y==�jOBy�A�ѥ��Jb�r�'�q�E��oR���5>ճte�v�:���9�(�h��	���%�'ي��3IJF�#� �w����30f�rsP~� ����]]�/��T�WQ�b�1��ݎ�8=E��mC�z���96�gJh�q����&�W̍1�E�+W��m�it�Z��s�ۘ��CaW��x@WN?��:��x9X�c�b�J��t+#�Mi�ߵ1�7�r>�_N��`9�����=S�k�W��u����?Vֳ�i����݋�*�oC�g,7���UP=V����$q�� � p��>��#EH�*�C�G�������������ݕv��0���o�?�� � ������_��}��ێý$*�~��Sf#��;?�� ?���\_��Y���#�~���rI���]��� ���� �������������� mO1�/%Ut(-�#�� �n[�������PS����r�,�U6_�^`>�� ����� ���x��~���s��e�@���s�����2�Iw���0��z:�:��ݾ����z����h��.��]nء�{���HX�A��vTA����u
UIuB�U� 坹��,�~ʊ1�}�D�'��G���u�q�Y�}7��:~FO^��]����u��:��gi=	�7�U�[VLL�ӵ�Ď�����=DݧSٽ)�*k[�n>�����/P*:,��)��#%�.�hf��c��(v��Pֺ��X����ٝ?�P��_ f�̉$!H1O�������p���G�N��бm�Z~���;y�#�O���wɚ]"�m.���ɼ�d|��XN�cqY�(���N�4�j���5���u"�R8W����!��,\v�=�i��m^��<Ի~v̎�*��[���5�	ܰ+�߅�3޿*������?\� Y�F��NΫ��o��ܣ��<�N��WQ��_���@�:Fg�`={pˬ8�
˦i0�x���CBI_�i��ё�U�#DRA�tM=%|�m>��ʁ&�(�G�V��!$�2��;�����t?3:�Ll�(#l[���U�R�u���.��� p�̃6��CN�o��elL�\���.
��Pw�4�cK��m�tI�����g�3D\��r��ˮ2ʙ�v�j��&������ϡ�>Fv��j���*.8�J �3(�}=��SZ�P�Xy�lXebM��|��7=+	lv�HccFg�Y�g�1���:G8�\��ʙ��U��X�`�̀kj��#oĆb�s:�&ՍZ���Λ���˓��/�{��:Yv�䟌���2`ڳ�UreRМ��s�V3:i�rp�_��q�P�S����w���|��M�*^sV��U��y���E���ldm����,�Sd�5���k,�h���̅x�h�K���c2���%ˤ��.u-L�y�?2�&��8�H�ϻ �z�HqF3$bh�9Y�AJg��.>-I�i6�FYpu75���i�,������.h� �O�e`8>76u�����]؆��΍��xƗ�n�CP��rII��r#�!�:E.>�c/�.���%����r��}��xr���^'���錒�JУ�=�(�+%9pgY޳�-2@by 7V�eV2B4<R/)��v9�iّ53z� ��!Y� �Ac�F@�5�V�Zq�'*�I�\�T��P�˾�n%��q���dQ�wycc��Ai*3�
���]�)rvf0�����R���-��(���EQ?P���UPT���<NB� ��,��X�VDR��V���gp���K��x�6��T��1J�Ǫ��x��J� 2��;��Mb�zc(q�VV��O0{�Ep�!����F���J� �Q){���$*�6�.hc�Ŏ?�e,K�cH����i2)�6'ȼ��@�ʾ.{4��HoLeM�2Δ��\�.M"|E݃H������u��zc�p�0(�9�Ȳ+)UiM�P�Te��)ı<���+��g��fZx��0��dX�G-P�@;!�1���ǟ<:A�=�&m�&��?���ə@Z�0_*��Hʩg����0	�U�Ƿ 褮�y�� ,I��A��;�`�x�N��!�+z C=\���S�Ī��� '@ؿS�k������2�Uj	5�Cj	�EfD�6��s+�v�,?f�x�V���/�f	 ӟ���c�,��X
�w���b����b�ܺ��&y/�1��>o�#Tɹ	�I���M�T�������p����t*͊�g\t���,��6PY�*� f4G�2�2!5���*3��"����ߑXY�a�?�U,�$1�V��J�;��XmС&Dy8ɱ�Q�'�o�rX�?���U�K�x�ŉ�	�
1؆pIeP@f2Id�+$��V_
ǀ^lX���~@�	v(�(٘����1d��n��:I䥖��L� ��;o�)c*┙e��!եt@��|�g�R�v?p#��1�#��YG&�qjp�9(X���W��U�oL`ˤ�EWE�2j��q�;!f�f8��)� �\���C��&�����J�	$Oˉ�#B����#�U%wF1���J2p������H�wga���%Xɘ�A���<���,\>�b�\ 7�e;�|�0rdO���b��72U��٘�'�|��0�1���`��,�%V��j-SC�Y�[�T-�N�a�� b����D<�Fh�?�ƛ�`�B0tW )R�� �4d�d�>8�����8ͣ?�>�o�e�Ƽ}1�����H��yRtw�2�-8�E,����jΙ�@�Ǵ���e]�Q^[��/.[�� 
��S&NB˝���r��<X�}�Gϔ(ذb��
��1�x#%�&Y/ ����Vo BE���~��6���"�^ �VJ��L� S����]g3��唀���(,b��O.`x��ܰ����V~n�dd`�Y~����X��$,���M&�E��'*,MH�;@�1b~X�3f�P�*FEK���FD��v�m��`�KǁU�P'��:΋Y3p�8O��),v	��N�����w恶�:��kEj�S%˛(-ES� iVٽ1�͏��췍,���Sc��k�B'Õ8��r�$1��˔����m�ډ7IQ�hEL�G~,Ts�>���c�M�4L�@Ɛ/e�*L0�.7���H��Q�H��/���K �@R�?+V)���^sI*/*���ء
�U+H"��L���oĞjd?�� ��7]��4CJ�D��/���̞n�y�E�F����}��y1��o/<J�������2Hw3E� ��E�|H�Ͳofq+��'$���e� 
�<��G"oLd��4*<.�z��sĔ�3e�B���c�I-���.��ȑR~U�;yk)�^4y~���Z�f� ��t�wE]���<�Z�",��+77j:�j���<j����m��5�2#9�D$~h�*�F�	dJlU/�=�c���";Q�l�Z�Ѐ�ggTa*�Q���~�:2���bVR�q���<��)��]h�<�Bh��+#Rx����-J%��c��gk1U�L��V3��3�i���U���F�{3`�-���9��(�Q%݋m𭷦2�t*��T��Ql|o&eU�P��,�vu�_�La�JO�{�l���#���	W�y|��T���d��).�����b�"dBǉ�>e]�+��f1�"A�kb��E���ֵI�U7�����	g�p�9|M1������>�X�k�/��͏���1��%+Y��3N���&"K�ԕRI�:��Lcޤ+�q��QhhU%M2X�
=��('�m���1���<��&Ǳ��gIIJ���+�5i�ـ����>,e&(�%}����ڏ��R�wV��OI�(w;L9E�qO�Y]�eZ~g6s�|��ES�@�f��bʀ+#2SS�C����4�x���0�Z�o��df1ȕ��+\p�Jc�2GQA-*|�yvT���%�1��9:#M&��eJ��>�[�o3��&��M�����Ƭ�-Y�Ly���8^��*4�iʐ�@��(;�U�1�S_�L=T.=Y�+]�򮶼��d�ĺ�O$+�R��"�G1���ݚ�ּ�+�߅��\h��b��srsqɃ~N��ػ��Y��g9���7.yY9)�7�a�bH^y�^jp���g,��s:s�����X�uw{�y�=mSQL?�h�W)���������2bω>40�ڇ設6?��R�i'^KP�mDy4ڪpyr�ɣ,h�3��	��Y�0ܩ,c{)��5�j�ש�2���HjF�]9��N^C��,H�Y2���(�Ns�:��6<�&�al�V�5�>�t���1�R���RQ��]~�o����V�k��Z�"��Q��2O?��������-w#�n}T�*�Uz#�5.��?�Op0g�r���жm�IL���UQ)�n̈�NY��	��OlomF�:��۷{�dQ:?��N�­�y�>��G�29|�ok�æ�T�wP*&��5�G�N�����Rڔ�}��i(��p�1�f�j5���o�g�KOb�]['�2��T�K������_���Grp�����u�v���r6wP����ťjR%���[h���쬲"�8�"@���@#4/�]8�����tz�D�^hh�p�Q���Ex����^�pAu-��o����O���:��t��z�B�m���k\k�_P�S�1���������n0p匲�LQ�s�}�]R���jR�&a�M�zx�VFD�@X�4��bgb�2 ��ܿ���=$i��j�V���]P����k'��S�R>�1
q�1a�u����X��C����k�q���zO�{b4���t�GW�zPd�=����ƞ�]J��Ե+�8mjc��)�Rl��u_U�⩪m�Xڊ+T$���1�#��PO�{<��(`�Xps�ۓf�z�ߎ�m_����I�K*�Z��q`�1�����Id��tO��WK�u�Qˤ� @�T�.5�v.���]WA���M	"�e���z�N�5�tJo���0�pK<A���{�/ 3J䟾i.���VU� v	ܨG"S�y�_�?A`���9'0'O����~���w�j�:y]m�����
h��������æNv��7��/�
S���L#4���ޕ�M��;57<?�J�ը�O�/w!��e�(,���$b��z��MŧCklH�1�4��� �2���T�d���Z1����;i���w��3�{�mb>޲�mC/��.�u�K�}��64E� O��?MgН<�P#:�x�X��"�>-������S��S�#'墂m1�C���\��� �*\U�P�&�v6o^۹Ѧ��T�V�<���iI�䕥�Y^#�tb�p{�'�=�Ξr�����#3��wD`����;bd`�u�����ńg���RM]�'3\�3��<k��������B�`��_�i`)��C�	�
��ڿQ��;�(M�,z_s�sN!(�ǘ՗�o�ʄ�/��Ka�g^����g;�u�m,WNL\�jY�iQm�=[W�6�����$�7�Įs^�j�5��#/$�3�#�/��<���*�G ���z�h^v�݌+�gk�9<H�^�ǶW�L'0�;���ކ�NW��h}�t�E�DԻ;�]u�v�E������nR�
��
a�x�X	�C�+�i����d�Z����m��R�k悥�JIf��ϒV�9Rd1�kH�@�߻>Vh���[�`if��+�X4v��wLqx�r��ѕp]^1$r��9���z3�]������ެ^����e�Z&��u>/o:~	�=����� ��2����(|�u{.�3CY��^����cv��t-�b��>	� �n��?[�}(�r���KW�Z֣`m�?-VD�Uj�-����,(d��*9�<rw8�gS����{u��,b�`��.��"�8�ִz�cש��8�g�QOG����gy4�bK^�	g<��uGX�;Д���EBTU�@����Ћ �}O���{�>�X��{U�Ot~�4�fw�� I:����S�t������Ϋ�5s-��nyɛӕL�^wl�-q�%Y���R�f����"V��lgKO�+M��B.�f�#`e�<QL�öz���)��yP��٦�*~׈�k4�׳\���E���7e%������A ���{�v������}W���=��ޕK��u��]9��>����Z�:�P��:���+��sȴ�e���?K�u�v<w���A�bx^*�4�E���H�=� vAk��v�}�ORv���K�L�+
Bf��lL(�:�H�֕��
P�]��w9N���ܝ?S�Nw�}E�j���ө��KW}7
��j��������㜇���0ڦI�����X�)�U�W���a��d��*������>��d[��;�6�{��EI$1�v�F6+���/r�J\��>5�I���i�ߘp�ҁjH�u�� �����#�^���?����}g��)�����>����R��q�rȷ�V2n;�i} tܨ�� ���l(��T「@�s�� ����`�G�� /�� Q� _�<��h�B�iQC��|��� ���z�C�'�� <��w����-�Vg�m��� ������$�����ߟ�z����阁q�Km�T�c�P�7�����P>��?�� ?�3���|�ǟ��e�=|s�
��n@�;#n� ~G�� �����?���>���ۓ��f����[1@U�x�� ��?������ϐ�?�;-�G�=��~���}��>��>���r��I�%�:Ez�V:M�f-3#5ruS��6m� �c�l��sx��>��G��K4?e$ZQ����/�̰��t�����c��s��oN�rí�tbY~N9c6�Gu�] �2�~VUfDs�U��;�ٯ�ۥ�s�}���}+����f:B�r�5g�ʜ�''�:�_εSX�l����(��ZT���vtw���]������5+�������l���ؑ�h��n;�v/�X�2+�[_]�z*�ޢ�]3I�h4�{��4`\�zB��3�X÷
�J�p�Kݗ��Ӿհ:��^���mc�u����S˞9�zB7�mB�:z��g"�����/"!��zM������I�F��~^�?�>y�o$��j� �� �4f��u��W� �Um����� �qPvs���xa�p-���Mx��!��w7�={�uս_��Zu`�j��nY}C2yHfp�o���A4Ƃ����!$�jZ��^ܗ�͙ ����4,q������>��zn�GH�:�֫'�rK;{i$v%�Ϲ%��G>ُ�=�J���I��_�i�FU�%K$ĆC.VJ�(�x5��VEcPH����Η����p�8��U�$�Y�5Jcf<�3�lB7����$���zc3�KhY1Ǔ�b�x�鑕�m�6�&ed���=g�(��	�2q�G"B �e}��Sg
yo�d�cd�uL��k[[5!u�Aj�����^kV�Ff3c�_�/9��'�������\<iҩ~s�Ը��ˈ��ۊ���f36t�Dq"y	,$�8�ƆL�U�WR��p����F_���%*l�ޒR�g��ڌhBx��,x���m>�2���+�
22� {c�I�^���˦t�T�o����J"cr�^YO�yL;���RB�.*�̕�i3Ɔ2�8����Db3���D���I�(N�IS�n���Țv��Fi�(����X�E�c�ҏc����p�$�6$rg���ejd4�M)p�e����8X��?�b�ݾ3s錾�&���>Si��+Z��P(���vg�ܪ�m�xŘޱZ(}�VvD��OZ���C�e
va��`���PFNP΢�J�m�g#���,T|m�ѹ!�7���������(j'�l_`�J�� p⁌4ͥw��FD-Uj� Eȯ!���P�w!�IY2&Գ�2����V��� ��$���~[}��J�p��y>S3��3oE/%+8RI	ȉ��e*X�d[��B����18�q!��K��B̛�lU��Lb4�ڋ%�>��q��Ku$�׍7I�@� �v'`��)7�Nl��9S%l�F٪'���Y� �u`	d�)��S2�I�8X����3HJr^A��Ld;c���I�X�t�eU�8�Z2nRU�<���f
XpT%�v0�����:R�������4�����F�)��Wc54���f�(�� �K�v{5ɚ�p�(T̏�:�|�QV��^����ѩDI�R
X&�^
[� �|�5�Vt��Yj(Ŝ,	�y(�lH}�T�m�H��r�04f.�8�i)J�x]ڴ�쎛��H!�D��7���+�ֲ���.3�RyrY�P�go�����ל�����dGv,�f�,J�U� �;U�c��U3��,\��ֈ�i�O�P">H���Hm�ȎC�eo�U��kg4o��[���u���Sd��͉b�Wf1��p|��/�����V41��Kĳ3>�_�4�zc$,�6d���*�m���W�7�� ��Lf-g��($�V�;*��,��4 �s�����`C-�'��$�%�6�҉�WeiqI�3ЊU��P�^;���*�~r.��1IcO�L���(C=8���e�?����)0�vW�OT-]�^I�!�Ѐ7o���;'4`�����1ި�w�	|��@��s�"��vD�&�5���6�N��V�m��a=�S���c
H��de(�q��1iX�u��r�Ƃs�@?$zc����T�D��j[f�4R�|SB��r�'�~��Yw<gz*�^2|�v�S�IĢ� ��Y�� q?�1�,V�kT}�:��+�G|v��=�͗�ʫ�n��c����u9U���T�DbEPv���G���M�ٌ=$fPY�v��AB�O��y���2��'-�0<!3J5|6
�I5���j��i�ꮄ��UK��735W+"���מ<otz��C�9��J�E'c� �H�W���P"���c�i��3��@*_�e
��:J���D�n�PXU�ъ6z�Q����\��C�l^H��δpM��)EQ���|6ş�ȹw#e,�1�gO jW�N�K�҉C\j�F���_��m����bk�
�.��ly؇��<2 �x��~�B� ��+������v��TF�4���&�,&w]��HP8|�L`�C���BlZ��>=vIǄ'/�v\�D�#pI.C8&2��F��%��\�T���,�71	�<�X��@Ld�[<��(��*M��ξFt�Y}b�y� nK�h����z�0XP3]'�^���T�+-���)j5g���,��FͺQ�N<�[�}�.� ·��2&H8�?�2"d�Ȝ|�n(���V,@U+���V )`�*�	��9�F&RjoJSz�Z����n~<~��ߔ�o��cד��S8�޳PU�89Y��ΥQ}1�y��^�
qݜ_ cX�/���B��]շ��,c���)p�#/4�~�?���6O��(
���6��c�%L')�q_ pY���|�	r�X�ʠ�c�}��Q)�1�F]xC�g4D�P�����9o��<���0��.�ڵ��,rDq��o)L���-fw�x��ȅB ��2�E<��P/:J;]Z�z�����ՙ I �������*�g,�|�V��5D2�qɗ��(`۱�H�`
J[Bo���3<���GO#;�3��6!��+-�%�ɦ��!q��-9����G �̷>KŶOLe	�j)�1�]Wd����jR��Vy�\��C���s��Ɓ21藡�FY�`؎�>C�����S��Ōt��3%	���h�^yx�� $���� )� �� ���?��b�-��q�!�m:-�l
�
�s+3�߃sv͟i��	�e�i��O��N�YJ��H��FhY�k%g�+i�9����i�o��Rh>����m@���#���,�� �Sj7����r=1���M����XK��&��G�0E2s_x�Y��&��0,b�ӆ6G���û3:���MT<v�i�q�� ���c��X[o�7$�QwdF�I�۫�%��B�
L�`���δ������A?/� �'q���wUʮ�s/�|LM0��翗����7������3ג�/z�:�o+N��4*��S�0Z���i��\>:�d,�L��h�95��S%R�����1�Ȓ)M�t�Ï�L��<~I�ޟi�@n<dCnK�ܱ��	��ι�_�\�+�Zεȫ0 ��L^���+��9�i:U�FVO2%dk(��!���K}9�������c�D,�;#�����|��Ο*�}�6� !���&<�Hd�%_UU�+�H�3ز��
�̴]�1�l�王�:R��q���&�ܫM5��+6!J�TS�i���'�oεл"���c��Q(r�L��g_���V3uOB�����0��,||� �S���R0P#XrD*f�U�*�3�,f�w?����eY�8�b��������mK_�5?��u�w���6zo�w˱����F���|Lj�'��cr�roF3�K�Y;3�\p$�4���Z��Z�M�٘�Ʈ%"�v�-������|�)�� �����Jr'��fo�t毃�����T���L�D�A�F+��hJ�Z`�'{���O�w��H��$d2�������Â�����s�]YC���2���e#�R#�gu;gޮ��O�7�2�����l-Z��9��|�1���K3F �Դ�nR�;�N�l�-WFz�~����_�
�~�����}��'Q��=��=R�[�w$W�^�Z]��f�C]K�*̠�Ч&��4���I��;��ǻݠuƙ�����1:�M�8�k�ex� ��n�����,I4A�ł�6�>�������������X�z�A�Ul� ���U$㖍�89Q�i�����+h{�D@O,\p���1�u���*��#򇦺�̬�Az��I�hW�P�~uu�G#��i%+Uo��$�?Z~ӆ�6�ͷF�:�����G�7��l���{�9e^G��U?H���Y�7F���)t�b��i�����r5���G�D|�G�G�՝k�l�C�� oݴ���ݕ�����N���+�]?����h�_<��IcK��.ژȹlh��|Lo������tI���R/�Y"���-��<��"�9#�2�*���'�=j�-N�ƹ���0�8͉U�E]'s�@��@;����e��w���S�.��t���辜���:w����۠��M��u,�;3	�A��?��cR1����^d�0n�uvn[^Z��WX�c�8-�}=wW-���o�z���=X��OA0�����K"OY�Gd$h��ʰ�p�,Aa܅@e�_#`be��WP�XYqeW��F��ssT�*K� ���m�
�+�R�^c+�xT�XrăǍOc�Ӟ�G#�Y�[k���pX��@�dQ���c��%�q��X�Vow4އ�2�Y�Գ1��uN��>HI���Ii��x9��CB�R�q��nZ�Ւ����ၜF�[H���8f^���+I�o���K�l��εVfG���A��;���c�A��W�S����#�����[�q�� L6����5�i]ßu�Ѻj�N��ek:�ok�d�2�j����Z�&T�Cd�"�q��5�b�5�1nM"��}�$Kkj��|�@LrE)�!'�㉬�;$qăi7���:�6ݹZ=F(�����I_�B�:f@T�f�"�H#��r��]>�S�GA]�ޡ�'.E'�y_���$�\CqA^�=�S��њ���}��X�;���<,�;�}�ےKrH瓚wz���%2�<F�����X�-��S���`�e����Ƀ���#���zR�^Y���E1R��''���?12H#'�H��3`�5��jmچ�'��~׬��5`�M�f����ߦ<	�����aR�%�H�JL���y� � �x=}��?y�����׺�����ܖ�m�׺���u1���zA�l�_/M���+�8��1�X�]=����gϨ���J۾� �,O�f�u�Ytߗi�Xڤ�%X�AVH^������#n�-���ڕ!��AdV�g�h����"�-*��{�&6"�!ހ��>���=���MG2�.���'K}CM�O�6cD_7�|9c�%6"�A*��5��-�Ǭ�$O"��!%T��g�-�=��Ρj���P�$I-�GR#��gwr$�p�,H
����c'�r��֫�V��luZ�t�S�R�I�.�#�]'�k9O�s2��:v���������(�mW��2��h����<���G�������#�)Ο?zY��i���Q�"8�)�T~y'��=��į��#��q{�нa��M�.Gv��:i�� ��-�j%���~&^�Ҹ�����G�/%[�;2edc��5�P�[җRhn��Mgf�-p���RFA��My��P%�٣�-DѨ"}�wN۟���ϖ��7��@FV����$��)0��T����lŏķp��+��M{^��:��G��꺕4�3G�;>��2N6��b�O�j��PŌq�6YMf�D��3�"��$ "�P?£�~��x� �r>��w�)�����_E��,�I�䷿y�}o�L=F/��??N�~;��wǭ/)�YQ�%��w��&�R��5P2�*G��TG s�����)�z�H�{�>����牌Q6bI]�����]���� ooT*�{�~���� ^���m+��2;0a�� �c���� _^��i?���ʟC�dYd�s�);͟�>��x�������^��o�9�Pw>������$fi�LX�� �S(��
�Fi�����A<����啸�
����3�H^9?�Ͼ㛹�;��R�{�����~���Z6�G�OT�C�~��~9ӳ�����˝ӽ/��䜳������AXS|�1�N�֟ni�Eߛ���d�Jv���걡n�4�Q������JI�K�#�C�^ޖ��������LD�X�Z�nض̜��V��4fC�߹n�tWi�u��k�f�xB�K�y�4]-#�)گo+$��yч�%��@R�'i���=�g�;i�����ٛN�2Ƃ$�)����9y���gbX��W�{����,>�ݶX
��A�:1vd��
d�0�k�9���n�n��h{���i�L=S��k��u>�\+��?��tג��U	ʪP�D�m_��imV�Og�6�+�ͫ��!	���AH�c���L���B���� �5�m�J)SL��$:?"E/�+&����?�ӏ��>g�õy��Z�Wq:s�4H���i�>e��Ej�yL]�r��&���;�Ҝ�!��ͻ�ı<�I>�'�$�d���g�g   � � � � ��=Y�{{�i`���H*b�w���Lc4�e��|(�;sR��Fz���_���K�]1��	c�8�O�fR���<�ܥ�ˎ���Zy9
��)�M�V3V3,t�K�S�fLza��5[�NzCI�ɤ1�!ZG͙/��ҔT�Y_����/�bi������������d�f�j�Grah�S�ߔ�~%FK1����J�yOӰq�Vyl�i����lZA���Ը�5��4S�Rr�3�:I�bVvŌ)�3gz>E4�C'*�∸�s�U��48�Iy���c3~�ғs)�����Ͳ*�mB�fRp�A�UJu���ːfũ$�Gf30�Z.d,����g��$\�5I�$c��>f��X�'�zc2&O�(���UfʆE�8O#VsPBb!��g�JNJ���#c=��U�y+Q6��� ����߆S���x6�E&ጿGNz�)�ⷞM\hR��@�[yk����m�]������3��N�5iLic�B������J�oB�\�r�/ ��r�匑�3��H���hƍVz��R����@G���qI4ܾKș��I4��.�$$T�8bq�δQ��CFif8���B�S'�����b�ǈ �,a�\pE(`�VU�9�y�MG�p����̫f��Lc+�3|�*�[��ދ�,���]�*��
��s��0�5�%��+g��9�h��k�t⎁Xxʻ@S��}�\�Ɂ��.,�4��� c����ٹ6���X��숫 ��� �J3K 2�*�<�b��n	M�o��1��0��#�v1>:�%�q�|�U�$��Z��;*��ޘų��1�n�TA4�Ô�7L�y<�7(���T/ٌ*<h�DK�BU2���5߉�R��/"�O�6`��Ujl�e����S��r-�����������L8ūsZ�&���eI1b,|d�M��6V`Y����VF.)e��J�oX��Jp���Ҍ���;��1����99 �|.7 <R�(����������"y3��w�b*�>#�0S:�����x�t����,{Z�5��Cʂtb'%|a����?��m�����9=�e���,�A�y2&��q���,��b�2�3���β+�}�xn�f�Uw�'��� O��q���b��|iC���T����*X���Ĳ��gBV�E��K(�f�|��U`�.�A ��_LaIf��j# Fu��+PgɏeR��rYIb	�2���Y�� %�"�g�vv\�� �?�zc<y��n�oGy���>~v
��l'�/-��n[m�1��>j诎��h��^��GP�?���v;���c	�-4�N�|tg�Ζ�"I�UR���
�!���KV^!��Vt;���*� ���܃��g%KQ��G&�2��yx����Ȗ!D����<'�b��N �y8!	�Z4W��	X�ޜ8��I����Fc#i�����-IQ
���]�1� ���)�-���:v}�z��ȦN����?���b(㒕EPYق��dnC����]րU����.UZ�`�F��( ��D�L�!W�!6��QI[�-
��~ .�);�Ldi�ѽ$`s��4ȋ��ɍ�r����1%P�7;/�"�
�L&;U'w��j��sȊ�� ��@Ř)㲄���t�y����WƑiM�荏{I�L�)�tām�b�u�=���w,f��++���bZ�Y�m�yQFŹ0c`���4��+�?,�C�*ҔV�1���<D�%P����㍗E�g��ey��0;%U������#�#`���f0�}�L� �Y�*�bůǛ9f�o
�wN\ّO��j�5�	ISò��YH�~3�41�s�� g �Le	p�|�7"��֥�����U��VM�^��9� �c$P���YXN,a�J�4���T���AW;n6�߰�%�Rl����^~B�\qP���q�n��4�}��� @F������e> �y//�[��S�>�*B��)7.ƈU˜�f@��
�PϾË�r�T�L�F�)�x���Ń�NfU�s��*A��<��trj�/�v�쪠D�#���w2~E7⼾��|1��Y2+*����T���YV�!���l�(�ߙ��JEM�.6fW�T_�X1��k�f
�f�,`�*X���C�x�S� �/WV�PUو]���a���)O#!��ʣ��#WĬ1�$XpyU?b��1c�ĭd(��e���pb�.v� �XĐ]� CF�ߴ�	4q��W�v��HQa�|�� �Y6B�;l��
����+z4J��xI	WR�s*n�~@�2�X�%_�bU�x�S��&�;�	컮�ȍ�PX1�x����q��kP�(K.;yN����;)x���ŪAo�g�*Z�o3Z�+D�j*�~��!<�R���
�@�&�&y���Z�f�T�h�Fv�||�ے�zc%w�	��%�ҳMh���K<���Y�!�_[��c!�)���iRg%!�V�PI�o@��h���;1�j�$���]f��g��k_�~!i�y�2m��� �Ei��4U�P��R�ʍ�6�;1�W&SP�G���a�uP�aɐ��@�`�S�cCS�\�\��G��y�)���''&lCg�\�z#�dZ��v�%z8~KJ��T�zO��E���&0O&����B���ٕ&]f��,�������j�+�4ϑ�+vG4�T,�A�6�����LdC"Ԥ�	�J���9*��H	S�/�:���Oȫ1��:N`(z)*j���R�7J+��NA��)<X��7����L�֗����������f^hR%A�yP�;�2L��K	Iʷ��S�-'�%�e�uI�l����JeM�Zդ����d�fG��+I9u��8�H�X�l�e���UZ�V�E#DD%>8�U��p�f�??�1�Rߒn�ueY<�#�V�ɢMy���%b[�9���C/62[2��fl L������8��x���a�� ��	��Я턓�¯^mXȷK�]��*�`�\�\���W��lAS�g@�m�M���k>��R�� s��@�jܣLQAWlgF���g|^K��xo�{r ۱�̑j����MeD�y�Tٌh/ ̈?�,wM��^��|ujQQ�Ɯ@y��,�eM���Q#��| >��i��'������/a i�0���O/ty3x
�_^,g��t|J*��2���U�j�YVs3�S�[1VUVڇc� 1�C�{g�e���#m�{�[aS��x��d�-�x��Rhh�-��X�j��ڶ���/3H��N�,qL$��+2������jK2K��j�!��0��s7������i����He��c�.���N$҄�,HvR� :5?�lf(�պ�HG��F7�үXQ�`�E*Q�Q@��
YGLe��=��[��Y.��Zk]3�����L��ˊ?/隆#Q�Z�H`F�F�m#\�tId�������ְ�� ~c�G�I�}���VY��Lנ�F�W%��'hmU��<�l�VX$��(�\}2��ʞ�{P�`4N�j�_Iw�x}�Ԝ4�Բ��^�˩�6�hF��(\�ꈬ�Q���>���'p׏HT��n)�	��4��E9�=��~ X-?���9�f�o��M�k��'�Z���G�X�佺�����r�=(�`�̕8�|���wz���%�ugCg� XеX�.�]^�8�N��q��	d��TޔUZPO�F�z���Q�n���%�j��w�E~��C:��&^	��,��G�{wH�6խ�v=�+In��7�O���Y�S���_,`<G�"1��}1�/���ӟ�۫�����t��rr_'
�L����N&V2���&m�N9�žM�M�goȚΕ^WE�=Hl���W �d wE G��3����5�dۺĒi:��r��y�q���x�3������8c�׼n��9��'Iv���?Q�C��=Ժ���Ժ֫�dix�V�TT��)�k�V1Ԑ�s��ug�[�m�z�f���n@�D��
�g�*������!FyFN�H=ͻ�)�6��;r�gU�1A�?��c�ƨ��i�I��ţ=��������]B=���A��;�r;]�Z�l}C��
�UL*�cdj��^�L���-�C�Q�¨c:E�l�"�ƂX�ޯ$�&Wc#&2��#PoLqɄ:��S�ڍ����I�^H�y���¼��H�R��#<�^~��c���5��I��-�ru���r)�n#e���ihQ�^N��o���?̨�� o�F����'̴����s� �~��� <�����r����=W�߷��>�����w/V��,����\<��|n���S��������66�F�7]O���;�l|����6�U�:؟��)�U%hy����lx�8\0P�˱�жN�<��^��z���iִV'/ľK��}�l�����g���^�{���5�|����z��n���N��L�[/4�i��F���z�0B����s΋�k:-����w��i���%�a����*��H]�>.YY�U ��Rs몚�ҥ6���!d�وL,$�ԉ(�
�}�;8!Cp����p4��]?��~4���>^��LܵQ�ej��>�2��k?PX#��Ԏ�؅'�W�BLQ�*��n��#��'��kwmƂG�O"�!A*��� B�}wx��2>w#W�/x1;�����΢�ɞ�d�vV��'2��:V&���l��jAh�lˮNB�: ��Y���h:��25��VB�;��Y��$����5r�?lfU�,rM配��ƒ��=-�v8��@��LEH����#��e�/s�%�|������� x�����n�.�N�uGI�-��J�@����X�n���K�nj�ǅ��'�z�uۥ:�V.�_sQ�t�I��1G,S��˺v��s��|���"�\����lIP�\�a4ȼw~���8�vx�;y��/_�^���0}��u�+f駷�V�Ke`�jc�.^��6���S~��e��s@qܪ�	M��n���s����51r�uH�~��Щ!lJ[��Q�bI'���=O�-jm5"�a�F�#\0<s
�� @�>����8��n�����M;E:>���i���~^�[V�L��в����������rk{6�K�r��5�5�m$�ܐ�����s's�%.�p�<�hb �ܕP�3/˫��,�J@h���� ��� �F4����;aC���ʈ�:8�:�D�r臏�2d�Ŷ�$��[m��ά�|�YqܼiP���n�O�s���,t{��.H<���<�>޽,Ĉ�L��J�� �I��;������P�G������1�<��?���!al��O!�#B6��P��� �o�?���_�y s�8$*�?��e��c/;Xص}3
��$�Γ��b�IP�`W�8�'q�>�Z&��k��]3L�6�v�H���ُ�8����� �MKP��Ԗ��QԆ!�w`�?�@ ,O s��R�D�'t1��3R�l,\_;�qt]O������z�
G/X].����+�O���y5�����M�Ժ�RS�%��fߊx�H׃�M�M!����/d@F�8Kvn-Žh�Sb+���+����i+0�X+DXK*'>6���o1�B��P�|�+َ��{�ߎ�u/T��n�����G�����������;d���)����b��>��{RJ(�u�r�j����{V���1��gs4�i�� Kbg%�PX�'�r/}:״���͡h�ͻ7k�#�&ie)��mF���
Щ	bJ�V���|������t}s����G蛌�}#��EԢ��Fǎn�k5=FiŢ�|W٢�Ǜ�s����[O�n��VբG��#�a��=�^��A��I!�2�o�zf�otꮺ��ԃ	n2p��bI���ܚՇ<3rg��i��#]]һm|��p�P���#� ���b�ii����w%����o�u�=���%���LK�w���aa��i�Ǻ��̞�Z ��
�j����B�⿇�O	���-��Y�11KҐ��ҿ��Z%	Z���@�g���hq��	�n���ɩ�dދ�Yk��#	���Z]�N*�������MFң�d�mI�lȬiI���& ���4x��d���FR�� c3���4عv�����Ҵ�N&i_�t�VSyyI��E7�By4z-��M��.�除�/��8��w�����԰�<&~�*ֺ��CQ�Wm�0��:w����23$���lv�	f�`4�f��d��qAŚ��&3+i�[�,yɼq��?7+o
&i�k5��׃�z����e>0�fFҴ��VX���i;.;N���i{5��5$B΍O�g�*��q���y�+<[T˅��*/js�G��=���;lJL1��X����!�1^t�E��%$+�8�ࢤ�)�/�>���/��ZtȡeFv������G5/͗�%B�˱�1G �)f쟈(��n��gj2U]�a���`�LP��[5<�:㜈cc!X�ZRa��������.!A,d�'F���Y�4�$��+e+��ȍBYx�X����S�XFdF��0j5��l�G�w�r`�|�UP1����&�6�K*&Aq���G2�4��O���m�i�4蓁�l�כ\,��j*�iUeVuv.B�� � ;/4W��T�VmJx�%L��@�0�"8"�Шf`�K�6���J��"ߏC���$��23|�]Ý��A�0�2O!�U$^`��4��6�E,Ê��N������ t�KV��Y��.��4�̰�;��C�G�(px����JqA��q�bL�B��+9���se�oͩ�pH
��G�I1ŚL�~"=<`�()#T���S�����t193q�M̑<h��zFK�,��#f���q�XǊ��
$�
�89�㺬�<f��Uظm��Fh��ec�2�,�,�p�Y�#"כ�P�	��g��@ۏLdL�(��F���g'YX�ʈQ�#��r6�q�0����Y؆�_6@iIf)_ɡb�������y!��Q�6�X:��(##4V�u,�i�U��3�gG-�c)��,)�ٚ�Z�,�"i
X�d�
��31�Nۖ<��,��p�հ���`��`�Q�_#d,��f*̛1��^Y)���a�#�7�3�G%��G���/�1*��`�_P�(�ȳA�.���fU_����#$�Ǒ��i��8�&ZNy%U�L[� ��ܷ$l�H�]�9��Ǌ"��ݛ� �x>��� >��n����`�X�x�X�gibȥhѹlW��zc���)D�c㬃ZtfZI��ƊM$	����0�,sn�����i����m� �����ܱ�lo�҄oiUj�y����u���~���A�=1��L�I�R�rk^9t�5(���e��h���Gbı�~�l�@�e&��
��!�|�&�N�\��B���0�*���$���xްw���3��e���j7dvoLa �r��C2	�k���R�i/����ąA�`���� \\d?���|.�*���w�ނ���-Y�؅�ٶecʕ�*p��	6�U
8��P��~����O���-�3�)����DT��c;�n��1�fAm�n�QF��Ŋ�јx�Ńr�L���6��PMB"�K���+Ld���T��nh��b`�2�4x����@����2��$$��<v�v4%� 	Cɕ��݀jś�l�ƀ�9�]i�f�q��B��D,�G�8E��Lc���3�fM�f�vy�~r�1���E��B�ڛ90t0���9�ҼaKW��Fgi�,�(0S`?��Q�oLc����&��2(#�CVd:����ύ��_�Hc(�Y�b퓰b�5ǎM�rd�<�!�r��pl �p��f�����D��IW�22�T�
ǼE%E8�Q]yM�U���M�[�EX( %�07Ɍl���|�i��,��VU,�m�b��TC|�f1`�o�U�s
�������PչU�gB�<?�"�q��)��k�QQ��ѐҕ� ���C7�z��p�����XmSN7�%+h���qP���`�vٌƲ�M�q���6���!��^s�+�⤒�(vY�MXə��G�H��Β�4aP�#�������(�0w�~$�8Ւ�5E$ʇ�y���1O �l[y����' �(�
�4+��$қ��C��C�@�܁%�p��Z�[ri�VS�RѼ�bg[n�7s��p7��_���JHd�r�_���F/9��'����Ǐ�1�\����!����r��\��J��
?��9��:;������+H�� j��s�6^;*�쾘Åg$(�,��Ƥ�ʳ���_���yp$�sRǁc���틑;ђE��yA(�r�$�O%� !��`P�$U{����e���!���)��tWnmA��1�N��:n��T�$�⢽��k��|���Y����	c$�s�kb��7�<�DUK4,�+r�w'ufa���D���3��mw���p�q��e��o��d��-lT��FiZ�F5)?��;*��K�]���� �zcI��<��ƴ�F��E+�+��2)1�>� ��H��8��|
	�)N%��|�S�x+����Q~��Aߗ�2���DC!x
5�C1(A/)�O��nT��3�;�ХCZ�'v�¹�I�E�F<P[���
�b�W�c+#�$��"b̭�d<�QMw���T�f���Y��OT~�B%̆��\Fw��E1؝��(�	 8nn~��2�?��p��x�Ad��b��9�S���'nD��G�dV�fd�'Ge�N� �vn r�+0���,���3F�=A����q�8�?�K1ȳs.Yw �@Q ��o%2/�<\_	�	˚�y��O�X������AR&뇒�^�L�^SF�Nf����2	!�r��c���<��e��ĕ]哰+��1� 7!�^�	Qq�tA����e�'�>B  �*��X�2�6f�~j�2���d�'$P�[��g�]�@� �#��a�����e��	��qUw?G<�9��fbcxsY>+�Y��q�M����@��ꌭF`9W��U吂�,v�u�UӒ��U�>�/m�r��( �!���z5D�Ӆ1�%�ǌ�c&�[����)PIT�?-�ȗg���l�m��&wbJ��lC����/"�e�3ա)�FM-�~�<�d�w	S�
E6�J��c,9�BRDʖ�����5(�U/8�+o�+���ȒJLg���>��,Մ䋑p�y�kc�l!9��!A]�,Ϻc5;�;�kBn�Е�f�xvŜs�ͯ[fdb:F��PF�t��F-�ʠc9���k�釙�h�s$�Գ�p�f�~>ݹǵp�sG��Pn��g(��ڍw�'6��k<[��m-�)���l�j�bt߃~3����c0��b�Ӥ20bj��������3*] ���AF'c�1/�#�q� �Df��9�U���R����{���(��M{*�y7��/���-��+��h.�B��i�B��w�G�!��ǨԍO��p�Z$畭dI�F`���}� mGQٺ��O[�{�~؄�u�H��QZF�5��D�i��?P~�}�v��޽�:�F�jG��3k����K��<9���S�P�I�H���5�SOm�wp�}e�5#Qax��^	���a_���� ��������Խ��v��ӛ��]n'N�G��b�긂�_��>��&�zz�oSH���6���\<Y�c�c�(Uu�g���&�V)@ri�!J�_N���Q̕����k�Y�n��I�V������$��'��g]��ާ4����c�n��ݜ�����<c�Y��Γ�Kw�^���:�3�z]�2r��k#|��j��,�3�6Nesb����$Skj�O��˥���+*�cS̑�߼?2R������g���i�ZڝMD�wi ƒz{��y$�*��p8#9ǫ~�}���;%����O��o����fN���!��֘����yz+.�����4�Y��s_Za��PA���Z�lR�40<��f�ZY��Vj���3�j��*1�^�	���'�IfΫF=�4�3�c"��Q8� w1���ƿl����l��;N��gU���sVڍҘ+�m� ��Qi�D�˜M9:���m��Ђ�-)&� I�F���}}��pn��x�x��]fC�^E�΂B��*��R ��'�������A�^���i�^��~.N���|�S:����ȼ�*���b1h`H́�Yb�}2���i�Mn�ؠ�eR@-�����?9M[P����~�Yו-�8'��۟���u�7��n��3�]��㋋�gQ�};A�:v� R�-����#^���iy(�bc���(���y���[���G��4� �
����K�Es-)�u�ĮL&(������	����w�u���n��$� q,5����vTG��p� �H��~���7c�㑬tj;��]#��~��~�޷�>u�\� �J[(b[�pꙀ*5����	]�����M5��֍�)�RUa����/^I;{���[��Ǳ�x�QInu���~��َ�ż*Yx�����{����^K� �Ys�t��|�KK�7R�'�t]���`�c�N6e��QWvT.�	� �O~�"h'��V�O��+��'� ���#>�*?��1�:В)X�j<��fc��� {�/��}�����/���o�}u�/b�4\��z7���{V�f��N����?*��Ȯ�2SP�G�&4WI���:��ke�-*i�ޅv�[vc!�DY"4�'p>$�Ҫ���D��B�t��}&���W^��l-��+�r�J���E��X��Y�qp��<��H�4�ұ�e��iyZ�V^�I�&����kS�Ք3'7B�R��Y6�p2Hm����<lZs��}��ӏ����>�,��1i��ԭ�/d����v�Jy��#����� �>Q����/��1���1��-G5��	ß����� >�*H�YdFR[�������� �n�]pQ����}�����Q��7�U�XM����.�$�?��'��Gߏ�� ^���s����>�a�5پ���5̽'�>����&6��k�ީ����:퍤�����S����n�����dlI�!2���w��*i��cPy�	$�|�T�'�h�hb���� f����^�zڣf�G�t��_��~�x2J��/p^��F
v#�7j�N�tZv�}ڝk����ec��m4�W��~��X�n���й��e�KQ���ɆkO �o�e5�؝4�O���g�w����$�؏�,B��f%>�Gb�U���qѽ����b�ͷ�=�Uz*$�*��f,ȶjz�L��4ѳFc�s�����ڎ����ڞ��Ӻ��+�bC�t��:B	�!׫��4�Y�
c�����*(5�O�gijַ^��jz���ס<��3��H�zC�����<���UA�6�-}���[DӴ
� ��C|�G�54��=���٫��i$>#��KY�r5.���:��w�Дk��tm��k��i�h86��<|fAZ��&����>��N�����>be�"����("_�4�>�?T��I����z���H�)
�����L�ؔ� �fo�i[�cڃ�Q Q�s����ύ�]��wVÛ��"{�+t�'�T��͏fG�s��4R�2�(��"9ٹ8���'�8���_7%%U�J$2�jwtٌ�Z/J��2o���}�,�[~>Dq���L-F|�w`���kSŌ�^��!���M-���2��|lJ�� ��T�3fd���O�/5�C3I�c3OL���Ne2�܍>s�R=�++W������,=6�a��O˲���=h�O5�[�����=�z�u�l}A3�c�|�L3�{��͎&6��JL��(1��=�����3a�^���+�'���ǎ����hq4�z](���C�x|��']�d!�̱�t�d�ݤ��R��yN?�|QVȀ����Z�W�9�i}8zc2�/Nx��U����KP�*
P���n�*!�fg�^(�fG��qe����2���������|���(���N{�z<UZ3x2h����ѕR�kZT���S6Lg���	��$�T�ՠ����H��}���ŉی�1�%.�E1�R�2�5U�Q�+�᫊�x�
��X�`�S�61�R��4�*6*A��ۯ�,rT����T���c,�7��ND����j><J�F� g'y�n����|�c.A&k$kS�R�	BȜ��[r�0]����o)�l��-T~ۢ~@4.�Q�+�M��CɎ죟��c)��fJc��������I͞�
T�URBm5�� s���|�eIT
�4��_�Jm�)`�o�r�6��1�v3��(d}8���삢�Ah)�o"m��n�ep�@j��E)��?��:�B�,��,9���f0l�`'��m�6�J
E�V�U��}غ�~B0��%X�yӉ�:��L!%��)�Jo�ũ�Բ�i�!UA��;�
��������P1�"-�< ��&@n&�H��3�/��,<g��"0*�1��cҳ?��ZxT�(�FJ�<���T�����i��X�+�.aeơ��4���R�.Qydl��1n,r<_oLeDdk��M^j����V�[��W!�wQ��x�r`˚4*�2E�����䢐,�ơ���NĻ � ���Y,_�%���D��KT�T/ ��˖�u��"�O�tX�51�*�EFpn,�� F��
V��]��� �0�Lw�g8�S�q�ң*����^-�T;��n�>��c5e�d��~ �ei�U9��}��+�7PP�ȑ�1�\4�Sr^,�Z�W�����@��;��v⡘�'����XK-�U�_b�R����G�.�x��mr����̠EEX���om�����EJq�U;E�4�f0�J��|�J�g*�9 Qf��)������&���qa������~[�l[s�w%~N���i�d[������G)��{d�E�ho��*��A�8��+��j1f�v�	�"���	 ~���O��1�;��D7��2��1f�ΛN�~��1gr�lėFf0�IxQ��!e�:V���B�i��Oo�`o�cԋ�K&W��&�6YE2�<r�&�1�Y�U
F���UV1�E��Ya�o�u3�P�]�B��ۈ4,��6ݛf0ԜMH�j�6S���*ʻՏ8��`���w�c�4��52UI��Z-�*�1i!#q��f?PIc��o;(�9?
�� �)|̝�0Ev ����`��5��i�:�TX�R,o�c���B�ۅefQ�1�2�jC�h�V�y|��9"�V�r�C�+∣`���8S%q�.Hs��D�e��- �h�����k� (�	`�K"�D�ڦ&o'�Wm�d��Yl\@�r�̿��Nn�r��fz�Tw��e��')�+����C�|���/�O�	��0x�ik�A����C�8��	ރ�K_�`�{�������(�G�9kG��ݾ�9�^E��ٛd�h�1�Ȇ4�J�ɐM��^h���;r����(��S��hlK
R�gK����+����'oLbs#!��?��<�.VwQY�52
����~J�  �Ōt"6/O�.@�~�fs*�����5g��^A���cq{�-��Vf�fY��^*�E^k����vnl�ˇ�dVOg��n��z���C�D�*�����5b�X��ʐ@X�;�՜�-e�bҶ�P����o�O��Li0�H�q��.S
�(*0uf,7{������F8��\1��`Yj��;IJ�Ie%8�� X��ʿ���h�I������fD,�K�D�� b�ubF����g޾\w�f�&;'?*1���$���]������:�Q�)�<|�5�@�@���(�k�b���J�s��ItZ�ך�d"+
V��w���Le��7��ʣ�ܨ,doc��㲋,�93��W{���B�*~w^@,��iJd!�2��� O�@��[����
�a�rf�<q��m(��s�lqJUX��~rX��A#V�:Z��#&����y~MK1A'-)�
&xc�2=1�� �^P�z��˞�$��1,��rEfo����2���h1���v��*���˛Q�c�~��`�n��r�>Ó�Þ^D������JЭ���HX�ήq����X�Q�?��Q?86�)ȰBܕ��d�e�����,�FZ��dO|�H����)���4g�!��Sv1օ(�M�ʰ�0��dY�#*2�T�"�~{pcLƮ��Z�y��'6'�&y�.?)%�1ݏر�I����g~ M����������T(IpF�),b�8p�*�l��@V*��O,o����pb f܉�fc��ѥE��`��{о� LIV+�������2�3�?!A���Ժ���'$���P��*�ds����5���6�QPFG��Ņ"��r�d���c�-�VRȩL|��>(����$�R���Iܐ�c߆�͢�!���|���q2�g@vپ0  1��LL	�W��Nj�e�"�c�����g�ɿ-ª���`��e��&��D�W<U�DG�ɷۏ���.��@k�"����'���$�D<~x�@	�,c#P]��Y��*� x��YhY��p�����l���12��̤�������;M��������O��K�Le�S�G�t�R����I���2w�M��錅uB^l��#r����)y#>NZ���Z2z.�K(%X���H[f�^W24D��$p�go]��pY��;0ܱ�K���Ƈ�)Z	ׂ+7=�U;���,ز�B�0tVW�] {X^I��eg?�8�ڈK�Iˍ"&�� 1��Q�5���E`�iIV��j0��,�6#��1a�ͦ2���Lp�RU,�Zt��nb�yP0W+�rAc!>��͙-�	Kx�n�eF�b��i'I�&m�`�)��l��Q�2��c$��$�z��8�+}O���TS��X���Ua8���s�WN��y=_f&�Eߏ
��(X�n�Ӂ�5q��ƭ�^��ئ���$)M��������-�]��n���5q*����Y!��!��sc*������"�o��s���05�;*ci��>��"_�"˖=��\�2&C�}iH�nF�X�5w���n�l�K2r2���>66Rd">j5�Y����v�����~f�W�5��ԧ<�X�
l��}��qZE��a�P�)������-{�:�K�ހյ���+7L����3Q�ȋ+D���x1�`Q�!��(Z�;S�4�q��.IF�`����$q�d��������(5=/N�iK�j���(��h�P�������B���4n���{b�quή��>�{���F��\����ö4u%����3�����L�ȗbV|�z�6>�����c^������٭�4��z?1Xw,I'����*9ȃ|h�FҴI��i� �Z$*H��~ր/��;�ڷ� (�َ�Bٝ�����O߭r��ݯ�M?+G�L�㉥k_���卓	��qr�'ƭ�-Q�}�ϩ��hr��5M1um:�]�%�p�؎^��/�3 ���=�)��_�ut������G֨Mⲱ��b��y�e{ג�� ��B�i��C���h�A�՝0�3C���NfWKh��Q�%*+^���(*	�m����Ǩ�K����^���4��n�![��sjD�����8����u>�E�z��4	��ۃT�O5��AF�� ���n=�D��g�fAꮰ��v��}��gK�N�����-*=;���77?3R��1��Ѫ$�����V0����GD�����H4O<�JZeOs]�$���h�!�=�[��Oj����?Q�h`W�mB虻�}Iu�,Dc�ߴz@����6bOi��=�cZ�^���K�v�R�'�Y}5��vm�e\��0tl��pq�C�FN���gYd,��8�0����U�O٧v8>m"�*Z�n��'�9T,�7Ԥ�Gܣ�����Ѩ����W�x���
֞	����%%_��C]�Ӄ��8}��O���&{ca=�`�c����F;�ƔH선�@R ���h%�٨*���'�?WiQ��x�s[�V���5(�����W����9 6E��q�}VS��ڻ-5�G5q��3`���V����&<��A]���Ρ�h#�]}��^��z-��� |p�}�e�?U��bP#o�F v���PX����s�[N���j]O��g�3�?Ф.4^���c�q]	�8���� �E���H�N|��!�޽�������n|���m����#����;r>�s�=��|얥������ѬC����L�`�Q��=f�~�Z�t�;���;���GVյ������]�����`�e2�t������ia�fKP������~��6���.���2�ϱ��iWR1F��xwN��D��R��#��/���3kZ���ODI��J
�4Qa�#�O#сp��x<���!�;+�>�������>�^�h:Ezs�}%\n��9��F�Ύ�4jdftx�"�ε���!m�lk_�V��:�;>=���,��[AY� ��KL�Z� 0/!v �h�����75	�z��{�*š	v�Q�қ4�������b��՜��&��b���?�qo����y��_ɮ>$��y���~6V��|D5uJ���k|���B�9+���~މ�	�^zV9���T����p��������f��Y�cu7E׫�o������rt��l�73�PPo��:�wM����!1���VX���{��H�����u�hm큣�a��*��yx�����9$�I�'�v�=N�d{�[~�?����|�IP�$]��f�Z7����$I$�9�9��f���w\u�y{U�N�hˉ����9�}c��LN�KCƆ�=����u8��V�ű�� �<<��yo��S@��9�m�kB��G4�UJ��~�����*���w�7g����{o閬^�P�
���7�;�GMt@�%(,�I�Fuow���{��^��b��V��Lv^��b�P���]Wˇ'��I���[q��h_|������������4X��`�w7g�N���^����R�&��?�#a�bf���E�����s�����I�c��Q(C��֕9��'h���� �u��y��[/Q�r��~����l��ӗ�<��z;�:���,���6�ر=��jw�f��I���䳻����?�ɺ!�5�B��WP���G(�Q@UU�� ~���)�fx���YdZ�@֘A�,�e`$�b��e�+ܬ����(~l��s�6GI���̘��L2�e����f�za�"6S>��RȩL� |	��t�\T̴B��/�ڻ����)���GI^�؈��
�z��w�����];�kQ�WÞq��U�Ī���`���]m����kAh�Gϸ�HT�35t�Ed`�N���l=6�-A����l}O6iE�a,��sUGb��U�͈�z�IbƦz^���D�p��i��D�1,~W-�4jVnw`K��k��zs���O�6Q����T���;�b���.�9:���;�4�9��e&l����kR��ĂV����T[4w�.ܹ���=(�x�f��%������"Ӽ�U�ѵ&��2���'�3��h� 2��+����>8r��JO�	ڕ��̼�����t̅-?+Ф��+M,F�)���>M�
"�_��y�)��p�iP�@�>H��$�]FS2�/��r�
quP��ɸҎ�� &`
���L+�"X)��gnQ�ؕ��㥢h��������~,�
�rM&��`�<�*8�+'����vSY��ΒJ�'B���3R9reخ���r��c��?�ŝXJ��*}� r|_ ��錦���e3�>Be7�RG�2��4ڑ񒢮O�jucv#���h��Q�v�S9�
�X��1R}1����T&�q��<j(�T��1�M ���>!��@J2 �����(�0<��q�dPl��9�`�#r���V��U������NS~L�=����g�1Ž1�2eJV�t��~Q�� b2��#O�?gZS�-�c$78-JNI�����I/*n�,�x�r���$0S�ڮԷ��n�7�
���R�@	���o� �cm�D���d�O*x�2_�@%�I�����b�V1&��q�s�<�f�7�AQrk� ���rT����|�����Ŧ�)4a7��8-/2���A�㔀�`8��W���5��1�L��f�H(�L���><��Ƞ�"�r.ܩ6�8�vX2�x��;��Q꥕����d~4Ry��y�3x�B�y��(�^ȴ�PWo�N౅jq<�<,�bJ�Y��-��mг��e"��.�۱�d���Vd3�n�h�$��M����7b�~�@��$&Zd�$m�z���0Q6�N<�F�Mx�W��� ��b6>�M���gX��&��s��b������cˉ
}1�J�y�"��bᝁj!�d%@����n�r@��<��[+��E����'%1���,��l\���r,`&Ч��g���f��H�҉���d��۳��f0��Ƽ� �k�6��+y
qD2�!���#c�U��"�6c�9ET�ՙPR��.B7WO��J�G�~�?�Lf2���Y��gF���pZ���j-�خ����I`� �!�9?��;]&��iX����� ,�B�V;1�q�Օ!��W"����G�RX������!,T� ��'�(l�!O
#&�r;x�)>8�����-�<}1����'F3��-)v(������*6��1��1W6e��M�r�Q3EAB�Ò��7~d�%�IIx�Ө�)uJ���kVy4� �tO�-�V0�a�f�%E��GƵ��Ǜ4�r����sO#� �Ĥ*��DSa^M��Tؘ#,0�\�*�YYK�Udc�cWLғK����YG�dF� ٙ�y� _Ld��,�VwP��N�(�
�T����ع#�)C�M8*�&�� I'��*EZnY�Dc�h)6,���Iy\M��!H|���dr�15pY�f��r*N%_�,a����㳸k�x��@U���,v;6��ƹ�=9�H���ub��fX�h�.F�?�N��Iv��ڈ|^:�`���`�QI�����c��y|1�a�I�ɼq��e͛���jŔ+�\�vb�Hc��,����3;����g���?.�S�"U��f0T�	��'z���Q�#�)��ZQ����e�89n�d�ք�1�d$��|u��,�9��]���S�g� ���1�+�w�R�EeZ��U��Wh !�.܉�>��r�2�&sC�qFq;I�Pӭ�ɳ*��&�Ɍt���f�D^�bg"[B��$g`���P� r��:�
�J��ژ��b\L�7��ϋm�*·�@�� *O�1�M�q�no���EW��G#�7]Ԣ����|1�ދ++�H5�*3M
��B���P ,�bw$�P�cJ�ۣ7
T=U]�3�8��%f |�cŘ�u��u��-T
�1�m��1W�}��F�M��z�|�N�N�gDuP�~��+�bP G�_�OϦ0�� Y���nʳe�1`Ri�B����iȒC���c�%��K�,yIe��f^u�R�pe��qT��ܹ�=1��-�gŦ5f��T���B ��g4"(���,x�1ʸ�dAFM�C3�1I��h��]������ ������v��q�r�� �AH��D�9�{VAġ�1����ee���M�pw�gH�`�u>=�m�G"�G�JH��?�)4�/Fb��*���h��B�nw��bXP��.�?�$��\R�W�?�̤�U� ���XǉM^�nL�w?�%J~��!����m� �/ �B��G��ݡ�eV,c�u^*�I�b�4��6RO/Lc�_g�$���1D(�DTw�8����Ö��1���e?��*�2j(<Э�2�
*��Bwr�@���0$�	��jO�q���dɃl�mD���4^;U�N<��݌v8�j�O�.�I�x���Ҕ|tM�s%������g�B���V	��.�˜�j7dR��x�ܯ�2G�2���pd���!�xI�k dP b���y0����y'���O�b��!f������.a�LeP������MA�N�[y�����v��C�i�0`�=��v�!n75&��K%G��wFb�ۓ��Y��Z�jc���H��q�K�V�9��m*��e`��� �Lb� U~r�Z�f� 4�q���#?�UBN2���e�Y��)�ܨ�M�|�%-?#�`��@ݨŀ�,e=Դ]l��0i��e`�&�J�M�[g9*��f0���)���i��"j+*1������U�A⠝�X�i,�3���\Nj�:�r�I��S��V�,N���Wt��#?��ș��H�㱩�S��sF�B=n,���Y0�x��IU�K%C˚v��,�@s�->sY�X�x|�Z�ѧ&�2��NW��&���;qd%X�Xȉ4]"������w�
LU���\����D�)�f1+851��Cc>6�61��C7�-����q�Q�f1	��),eݙ^TvT�FPU�;��?<B�2%�f��*�I�5d`���R�J�`���b���AT�F�����F_������6<Y/r������R�#^y*��V�NJ�MВGx�w��*aE��(21n��7�>��_s��w;(�$�=1��:OL�Ʃ|d�	�#8�/�U���9�M6?~a�s��c5�����N��c��Ѡ�G��vK����
�����NP�^3t��g%{��� )kg�b��l�yWi5�i�(���I5ur�0�rK���u^��\{���u�x�g�)��_���K/S�lX�9����$�~,���h����=w,(X��T�mǦ3g}���]��i��W�R��˶�� @k"��+�㳥��Ż�iY#��Yy�A�}d�^�F����]on�2|���r������sq�hO���h����}�SP��sO�&��	�u*������չ爬�4|��,�gҏb?T>�{��ӆ;��a������4�gHf��%�<��]b�-=����1}�v;CZ��Q�4�u��c��b1���D}�O�d�.}�V�-٥�{� n�>�,���QS.�ň�"����{�e�E�0�Ԅ�H~����?E�ZO��?V���������V��e_����Z�*��Uv�w�}��u�cwim3@d𤐺����Y�x���T!O���9;�?p�;r�������L+�+�8O�h���G(G޼�>��JW����~��Dtޫ�i�օ��T�5��?&x�&e(�\��wbCr�z�����u��
=:E�8�D�p��'�(~�O��{j=b�w 8@ǿ��[z���W"9>bie�]���t����D�{Va��C��~��4Kړ����4%-LLY>NN<�tz�p(H ��u�/�h��ļ�Q�
�B+�)n��ߦXtH���N	�ef�nO�v���=� }����Y�܆�ێ���۷@���V����y�j��=+�4��Z~�����G?UwD�Q4�zҽ��:z�����U�fğ[/�GH�T�{��Y^BO�B���{omR��I�j���֤1/Ҭ��!b��U}d� Ϝ���Z׿V龋��uWQk�y�_�k��,��2��@��N�����m7�W�w��y��#PB8A�5��Y�׵���Hё����]�$�+K�W��R7 *��̹���4Sp�b!
��+\ |�:���~�"�������wv:��gc���S�:w��F���&+�Z���4���J귫m�j��2clT�M�.�Rn��u[Z~�Jͳ��;IN�Jc~�9"�dB�F*����6E���B�z.�QU�Q4%��Z7������d�3/
W��~�1��u�u����ퟬ�>�`�Q_��CW辢�^��MZ�֝���Y��,�Aq�%]��x�n��z:04�χ���uC����ۊe��Id�%��
�ZY$�̲��"��.�]���d�z.��$������$0٧�!���Ed��D�L��7�Lй�ۏh~���ۼ��е�����.���9:A&��u�e���gU���L���<�KZ�L�z�m�,��|Q$Õ�֧'�}��/��n��5]��k֔AF��X&�3�G������(��/2yQ|����v��M���iˠo�$��U��is�#��a��а�L���s:��6hc��ri�n��:ơԙ2��s�n����Ͼ���֧ ���j�v�~~S0Y�"��T]ב����Խ�>��Y�ml�����f��0@��e���i���W������g���{wO�r�tIH���*��M<���F=�p�^ ��V%�p��{��֩���6��{g���p�\N����՚e�o���1��!�y���B�j�;*���W��Ι�(���ߔyH�����<��-�?-{� �y�/{#��������K���Ȋ9�*��U��&�y#��^� ��/��ݹMQ�LI���$���e4Ȱc�+'�j�>�jA�Ĭ_��lv���kNvoFN+f�"�.�d�-1����o+]}Ȕ�&HІ3d�[���4<��u�Ѡһ6-r&���,R8sb�P���wdf3/�(�0�ڏD����d��G�e�d�ho!���u�@��D�M6,fe鎚ˍ��-�WǞ����3H����Os"�<_��RV����C�A��L8�d�䪏�A�r�`0��LyJ�PLcB�(�#�Z>���2ɾHȆta�0Y�����R~)IN+��7Ph��c3��1��/ϕ��&|Ʀba��uF����;4�e�7�m�Gv3-hZ<!�1(��l��1��J4Jy��hQ��Y$�9��r�Y�̉��X��\H	��)M[#�6��)[H+�d�g��ʩ�J�W�X�O��,o|Ge�ʞ*�f��lPER�L���M��%9�X�a����턄Sΐ3�1i�W���!?b��#��/�_�,e�Brǝ)lI��j�E���b����7Ewcʌ�6$0m�˜1��I��@�F*݃�!><�
�����ۊ�
F�2l�!lT��a�*x�k<[<���aiy���n�wcĞLd��Q�1�JW�!yZb������Q����wUS�bwc����)�,�cc�4y�ۡ�1`�%�0��䥌���d� ��Q�VV����'������t�Բ��W�!� j�IX»H�?�:�k�URYUro�]�1���'��]�q<4�C��*��$r�����dj"up�I����B�Y9AV`�dU���E�[��Ǧ�
)0��iӐV�H� qfw q!���RX���\���F�J/�j7�ܰ�vf	��1X�UUh�?�	���K+�n��S�!bv^>�ʲ�D��2�6��z�j�&+�M�'
?�Ϧ1C���O��ϕFZߜ��8�)������0����֏G�q��Fr
K"��n*X�'�o��r��DǮ6E�XR�G�s��dfU��NoNj
qc=܍�� kx���|��|�Y3S�U .�)�l��/6P7uc*\��O��ɢ
�w+1�H�o�p��݋����hřI8ԛ��Ky_�U�ʳa�&��r����x��F�eY�r�
��{3S%�4�r�!��F�@��,d�3��[�ψ�Ê"п)�U^k�h��7#c���i�X�Uf����A���x���
�(�� $02�\�%P���ZlQ��eM��,�#�����X��Bn�C�B��[�.�PѓӚGɳ-��1�eٌX�sv���J"�utB)Ctm��T��A �Em�c�������
�;!t]�)c��i����zc����6F;��(�]�<2-J�	��Pǃ��sv��M˱�ũ��2���*��8���S`AR>���D\:�5Uq�UuH� �� ��t��$�J��	JeRᑨDG��YQNܾ�v�X�J�$��f+_0X����ڼ�r`U m��&�D���*%HDDݨ|��զ�%�&yqg]��*�� �0#��$|S%H��(m�B����r�y�X,�u�n�����v�&2t�/�+o%Q�$mJ����p��vn$���b?���ee��|��5`�fȃ��?M���!��+�	'&e�rT�.�TG�(���q�,�e`�$�l(,b�#�Li5ƕ���Vf�]�8��HI��W���V[����Onl�I*"��#�����C2��rM�����eo�V08�d�#>;B5/J�|H���g����U�[v��Ō>�����T���	��6Rא�#��%��x��6 ;D�6G�bR�:y7`O���|�����}��NY��y�X���+���"M�_��S�\1%x�"{ցωLc_)�;1
1�����ubU� ��M"�ꍏeu�U�G��"����Bp$�@N;nX�BB�	ݥ(���BG*�7f,�76g��T��-5Ph���o�����"���� �I�wrŌld��gV|����r�/��`�&·ʨaR^?��j�J���UR�&��h�`|�n`X��� M&�ʌUI$��E7d��G�AFr
��Y�)f23���"c����
 ��T	F	V�S�*n.ı���9����g����"�(�;�����oLa�Z��|�x�8��Q@����&X*��$[���錪:*cҼR@�H�i7W-��&y���t
>6* c���K,=�+l���ZV��l�h<I�>0K3��e<vc
�y�Å)"1�,��NM�Üq�|�<��a���.�)	-��U��Q2�$bI
93q91��3�w��TcΕ7U<f�
ń��n,�Ġ��4!��9��ڹ��d#����TP��s�O'>�Ɏ�gf���Y�$iDv�PYRD�f��� �$�*��R1!L{��H�Ū�z�ƨ�h�����?��  ���c|�2k5E}����ȴ�wY�Um�\�Ĥ���zc	zp�'3�^K+*GsW��Mf���y�ߏ��1��ڔ�%ނ[Y<�9�c��5ߓ8��^����9�3YͶP�W�(�dS i.W�e�r@f,X�f0�g��Q��1� ��4�ם&��(�U��1b� Pr,eJ,��E��?-(�%��1�rj��T$���<��$�I`�eP��a�Ep�Q�v�����0i<z�L��MG�5.(����QR��?B���.�T1���Nrw�ʵ(*�F���:5QC:��ݸ�8�4zc0�vR<���\\��	w0"H�C����Y�ݨ�\�h�޴���r^d��Y���5��X���F�ȡ�(�lp�*+��agI ` �v�X��E�c
ai2?&CR���zYɏ� <�#n��P����vTWu�J�J�h�W�I~K!Q�r7f}1�YQ\'�Q�y��sTT�&5zs��'����Nf�_���W�(8T0A�T(j�nEX�� �_�v21o$r��Β���Q����J�n��Sp[��bYX�I(�*Iޘ�B5��՘�s[�H"(��>3����Ʉ8���0D��9
���&�M�f� ,[��1㠤��	��Fn\.Ab���E;Ax�� ��c�-g6��g���>�w��rM��<�%�[�%�,��T(�b�Ǌ2P�~�F]��(�������c��+3&�El�,ai!X��&����|:'f1�1��zR�_�Wj��ZC��93+�A�ٓf!���ݝm,��F��O,��\�F�8*S����.�k���e'��W�*$�f?������l}1��(����J�<H�v�!������T A!���	f�2Rt�O��;����J����� {�����_��9��K8ƕ�l�T	��fu;rpQ	�����X�p��+GH�J� ~S\����e`F�e�,�+4�*��8ad�����f$��8���dc�W��j���b�m%QÕ�`v��*ys,�W�֌�a����R�-"M6F$SƤ14;��Lr�0g4���p� �ޡ������6ۈٛ�e���,�hd�Bf�8 !J���:y��EUT�P��?�����X�Z�x���p��Z��CG9)-�B�kGO �/Ȇ �c9��_jzn�JQ��_*�V�l��rH����6J�Rzљr"�~ip�rc9�?jW���Li�Z����MBP��Ӎ%[��En.Ɓxт3ͭw���>��\k��N>O,�(��ُ�$;�#�P�G�1ؙzf�p�->�zf���l]CNȶn%1�0�DZn,��3+�@,��@��y����={5�<rF�$GSʲ:�����H#�s�h!���B�+�R�G"���ÆGF]z*����쇳�ׯ�M�{S�T�/m�GB� �_���TϤ�:�������%�Nw��w.�^��yj�Q�UթW�<wjUԧ͒8��=�@_�,~0�k�2��zt�ͥ�vm��-@�f�d������Yh�ǴV�;m�� yY0���>��5/�"�F|5} e~��u�2U�ȻQL�E��q��ٳ�m��5���E��)@��r�N�{$R;e@G��uZ�w��[�tT㾴�`ϦC���]�ӡ�^)����}��� pA��Ht�X�~Z��;8MZ�/�b�ruiW�*F��ٵ��k����{��#8S�6L�q��������Ө��J��v��x$k0��;���z���%��~�f�{��gn=�v�/�p���>޻�-W�zs�]�����t��8.��隖L��~���c��Ƹ�%'�2q*Y�Iz���\݋Xҧ]?[����T\�5r��ꥣb��h�$�jҖxd*�F���:��G^JW+&���)$�^v��ʥR�Yӻ�eVe��H��h\+�� Ёw��~��}�t����j/���� ����sk\.�mOȫCS����o��U+4k�?E�x��x�;�=~Es��� ��3��3���pd#Y
�x*� ��(#��k>��w�:S�?�����{�߾�����XEҵ���.�n��n���]+P�����ȏG��6;f�L�̬�'��/2�1GJ���V��a����-ۆV�*��f�Ō�'ખd��;�)�D�~��ޘ�h�{4�������6nZ�2��r�*�D�bf���^�)���];��ug|�������]*�}�j:��v��_����#/M����K��8�ŭ\R���[~�W�;/�[A�Ne]V�׭1":4u�2Ia�:�jiK�,1�V��2�Y��v�� �^��uc~���{���Q"���7
�׎N�H�D�}�J$���w�7M{i®fG,�kۦ{��P�2S9��L�����*��u&KZm�_z��t
�俾n���j)�$a�V�oG�r֬��y�vĒ�+�GB�Mת�-_�U���Nb-��+=H$�T��z낽�#}<�O,* <�?������
u�_u&nUq2t�Oa_!4>��W�I���U�l��d�X��-op��LP,�MFc^�q�=�w?ښv� ��)i�;��44t�W�.���
,޲��X+��T� ��Xc�~\��N���Z������K2������dѡ��^ ��I��m�gc�z�e�3�I�>�V��Le�v��N�fM��9�)m�L�6.�O�J�,f��f���;i��t�Te��Y�`��yM;��%2���ۛ#U��]=�N�Xڂ�1��sᏧe���1a��g8W˝<z�I�TIR�NoŌ�]/�S��	ۆ�����T���gľ:�DZ���|�]�N]U c6�4L�����P�kRk����r�����q��f�p�P�e"���v%����o�����F6���l�o���Y��<\���@d_���Q@�X��t� ����<:����j�Vճ;�+`����8,��̷��R�?�y�.��B�Ԫɤ������h�5^cm��3"��[�:M[3�c�2x���L���x��Ѩ����L��z�����cZI�ς�c��k9��+$I��v ����g���<�E#f޾Mõ'Y1Lq�_�r�B %Wd��^p���;`�iK$�W�<G��@���g<� R�ٟf2b.0��q���!H�j�'u�C�C(R�9L��m���s9�Ļ��Ĩ��;&14���-���H�e�e�"I,��\)�� �X�B��o�,������	W%N߶���C)��#Ҵo ����7a&��A��������:��p��#4�Է:�����i�/�P��Rd�AT��.� ����u���HF��Գ��U�F�m�$����:����C�&a��Fwv��Ǜ���˶������n�2,����U7>d���^3bN�̃�U�j��xD������
O
��5,�󬛊��>��=1��(�U�)oˋ��(K���H��QY[��rIcAWVd�������9�C|�	BR�>X���*X�(U3T��,�\�K*I�@��UO�f`��#E����21�֓dv�E����M���e; �_c�zcO,�i�y���J2i�f��xSwp	'e�B8�������.>̻��ԉ�գ̅uKlP��o�<�T�����ZhF�_�x�d�Q���f��9}��.�`n�	�I8�O�D�(�Z�D���	�n8�j�V.���AEz�J�y)�����r9>G�U�J(Ub�,a�),f����4mpH�5!y}X�,��7�22*.0r�T�f���(T1��X��x(B8��r�v1�5��J�M��4�Z���(&(��T�o��!�G�LZE+@�D�n�)*��,I^?�+n�b���R�֋J�"��V��'SYf2R�����oLeRUEE8�:�s,����T��W�0�	bC���|�c�E���UL���n��h�7�yxl�^M�>ѝO�Y,���r-F�,*%%h����!r�l>O�B�>�����Z��"�//���L�.�ҨR#�-���}1�!�!#B9�Ԥ��S�G�#]�� v*T����L`�x�/��1�|���� ��=1���L��Z*�!��o�7�����e� ~���څ�K34yƾa9Ჷ�O	X��L I}�݀K��[1��2��Z�a~©s>TaV���b��Ԗ!�b�\�x��4�2-e>97��\��e���䡅F���1�ƶD������L-K��(1�a�eV~lx"���dR�_j�t�~Cs̜UK��v��lW�}B�����I�*�~V�*/>e�ߐQg�}ܩj=��o���G��vu�5�8��kH�9Cu
"Y�UBL`���笲2�X�D�r�W�}��m��S�m�l鎵�vU���܆C��&w�Q��8���ǚ�0�P�U����ҍ�vI���VHÂ }s�2���Z(��֤���#���rvi���M��'�|Zdd���m�l~S)%�8��Y��AY�����ʲׄ��r*�vt(��,F�x��<�o�q��I���᫵�ƌ�J>3(f"QNqgB̤#�O�2�-"��IL���fȴùj=F��'=���
~o͌s�Y�����q[��L���j�2�v�(��+���1���iy�q�,���+�U+�m�@��n�W���o��Y)j�E���U��D��|�_�W��A��GU�$kN	6M�L��-�@�YVQ�5� �"��Cp���M<B���mj�j��p~%�)�t ���AO c<���z�L��n�NԸ�_��UT,����ƌ�BG�@,�E�O����7Pv#t-錩����!�UH�)���LYJLrs�W�n@l�I���ЖzEP�������93y&WeY�f��lXȖt S��Y��`�j*M���<MP��q�%x�d���>ʑ@�X��c7�+�h�if4e�6%@Wc�6z�|�E$�iJ���d��KQ�vŘ�V)�k6&Y.�&I9�y0Z��a8o�؉�������`�Phg=����]�z�3��f�w,T�0��Fv��b��nY�y���ǣ���6~M�Ā�� '�ӁEXx�*�x���5��lSv ����V>��Y]�gLcr�-*:��v��IT<UJ��F�H,a&�/&� )BydZ�P�>fT�f� �d�,��ٌZ�#V�(��*hckE7ݘ�\����6�6Ž1�I�N͐�V�DZ���> _����������9�$,��E��r�k�ޕ&�O��?������� �I�.�	�7nIMk;�
���U<څ9�-�[�?`����t_ƙp��N<����xC? v,W����24Ҏܔ	�L��]��n�^�O#��wP]�&�zcq�F����[� �Yf�q����3��K20f#�Y�5�ħJs���Szq�%�
;L�i��W�����[���f�|p���M$���fnd����m���w߂�4H�aU�e�� '҇���U]�ryzc��8֮�j�ZT�gG��SI4kT@�e�UX.�O��hI��M���Ʊ�P�J��[���n,6��̑�5�&5C' !LѦ&�R�)������3|��*�Uȣ%���4Z�.o�VI�rP�vu'��[2��fðY���v\�u+̨���܃�ǈ�����qݯ�����ݘ��Hc�x��H+��,cLh�ˣ�h�Ԋy�ڪ�Ff��ʤ0
@�F��cн?e�M-A¼��!#�*�l��]� �La��j��/	R����e�4Vn�������Ē��Q	AB�"��0��>n㐡�n|�ǟ\HqĒ�����5�նu�`��ȉ�R ���p��`7��c�!�|�Zg�eg�Gv~B�ܷ��l�� ��c��Y���jIh�Ȯԡn5�N[;�� `��I$�0���SI��u(YU$kF`O.c��2��cj�Y�b�%�@.9������$���C9p�fz
rI��2�o9(�lZ��7��/]ԟ���c�EZ�O�ƿ+:91S��,�8���r��^�3�>:1�����C�Ȇ����#���Y���c��T(��է񉗳� X� y"��6S�,����
Nrg�Y*<l�VI���t%\P�WةB(���P��N��D�Sm@
�y~�挫5e��|&�3:L΃��͐��;�4�މ\o�&��<�;>�����M!IV�&5��z�"�,��;m�6�wR�x�O�0uI�s^J�~S�:?5�Bl'E�B�#/�lX�c5/������-�\A��Z+���RM�z,P�P˒<U�<]��OF3������됺n���Ӄdddi�v4Ė�t��譜��2
cᣀv,g!����Y�1�0�$���	s�>V7�U��(�����ES��=1���m)�U©L��Q%�D���eUa��O��Xq����ݾ�T�Y:�lz��2���]%Z�7������S�"�n�T�Tn�1ٻ�tl=@jsSz��﫱/V��R��?#�q�*}�E#0.���euCF:.���� ��^�v��~�Ӵ���ʩ1I�2�"�3�+���P{?����������[c�<-[(�ԭ��hڳ$�$ce[M�*���z���z��Ղ�f�ު�R��\`9CB���(#���Ѝ��5�e��_�y�5�$�ߦ��"ގ.o��&�J|����n�I�L�Bv}0tzz�F���:�z��	�_43`��JI�]�_@
�ԑ�b}D�N��VZ���Ȝ���,� ��?w!�pyf�n����M5=����'�ax<�~�Լ_s���>��-�O��	��L�̼�~3�J߈tA7��%�o�� o�>���%?�H�Z z�ĝ�����YG����|��9�F/�mU�?/�q�������ǲ=q��]��:�(�[ҳptkGT8z�>!Ѵ��e�YǮ0�6�B�Vy�;0ܟ^�����m����\NIVWW��=�ZfF�w�����O��.�mj-�n�r�&���*#G�e���n������?I��o�G��t���j���~X��-W��e���9��H�u]I7m��$�{;6���A��t�O��f�_���_~JzS�yY{I[6���h�a͇'�Yk;V� ]5*ֵ���UW����P�����Ӝz�K6�]"C�<M��_[����s���]�Ie&��jlڍ2r2ahI.X�!DB�U�W`��ڞ�~Ϋ�^�Q�n7t�Jŝ��}Ң�D_�(�'�F�v��KFд�t�'NA�ƱC¢���f<��,��I6>��.F����_�Ʀ_���q�k���8���*n���(T��
sQ�ߗ,�Ο�>x�8�P�/y��\�4w�\�M�pc�D�_������1��H��8x�L��4�q��zn'�>><湏�A���� �F�@Ns����1���<�`����3r�.6V�X@���p��Ft�gؤџk��щgy+��-�����65��-0��izG(6=�,˴h���Hό���f��F38��I>>B�|�Ƙ�cRwȆY��^V�9���bquU� �fc3��ӫ,�Ȝ0�s�-I��#2�L\5���d�v��(zs�'�M ������}=�T���HF�����#��ȱ�ĕg���� j�>� �1�?Kҙ��J�mF�ǳ\jR�zIk�y�B�������3��钣�d��M�s���:; ʛ��K'�S�%S��V,g���ZI�;q�|�Y�EaW_���a��G�91c/�x�j���b(vL�6��ݪ�U��A�ʬ� @��ג��_*��v�s�lu(���qb��h���&���p�C(f2`��yY;�!��
DV��Ѿ�R��r�HP���|m�4(��
�Z�=�J��T�jT����,x�ld�-�ό��?5Z��u��e�#����i�lAc+Q���x�g䏋�Lړ��
1�]�������>l�C�̂����J;�,ӨUbAS��Ld�x�i_���`�1>G�x�s����<[� Ϧ2+��Q�Y[���,��2����������zc���Ŭ�r�<yJ0uph��K�#fU�A��>��)�x�p�
R�P�dg"�����������Ɯ����jp�"*,�� NT�)�v�l8�<}1�%�U����'"0@���!AR� B�ܱ�����T��c+4�`�̛Q��7��E$�py��#�QY7A��)����YL�j�e��!$��`�1Z�8�)E�PL���=�>ב��"���O�2�7@�=�\��.ԤkV�NT�H�'��\wm�;/�8�d�Ld���vi�B��3g����#��~D�9]�}1��_1��,�*U��x�C�1��D�6ـn,97�&02|�UZc�ӂ�PZP"�I��j��w�
�	<�ر���^�����Z+��;	�B�⣰j)*9������ ?�TZd���r'#H�+A&f4�+ؤ�U�r6��$�N�)#��~3��l� ���@��ó�n��P�a#��'�Zڊ�i+R-PW%��g� 0
�,c��O�J�y��oD���IP�$����Q$g�')^�&!�&@F.y��V�|�����P�� r��PȒ 1�I9v.`?miO;����M�~�ŌJD��[�.��`��"��E�
�@GR"�v*�T1���P0&H�2-��2��i%��٭��?�'v��;�r&�t�[NY9i��
 �QX;3��>_�%�=1�^u�rQ��*X	���)FD;�8;+O����X�6���ʨU���4�N��n6�� �� ��᫄��pq�!�=k���d�h
Џ���\fQ�m�Y��$��PVV��'feF��E }Tr�| 8����bq�T��W����mY5�b��R�ly J�}1�ZR$'�21�dF�e�p#���/�/��rP�q�q�Ȣ�R�U~S�-�X�,���N.�P��g��D.˱��S��':�d�1ځ�,��2P�uƕiuX� �Hdx ��e�2�Pyl�����9��g�' �M\s��22M�<��;��X�ܶ�`�2�I-J��'<d�����迎h�s��m��➘��p���D�R�9 �Q�v1�C��QN���F�);�1l,�JN��|q2�E�����fb�YJ�vS���HF\��~�T��[��Qۓ��-ۂ�*?�$�LaL';P;�p�w���V2vkr�姙\0 !}�� �c��Q}��B�"�w�!��(�W�$�o�����H%����n�E�G�ׅ+Bƕm��F��>�f1�)��	�_*��

�)ƛ(}�X/��&ĉ���|��V��	�^E��re�o��=1���"�Ӧ++;��e���񛍕ۄO��l۱�}1�xr�PJ�M̝��w��m51���X�rb��	 /)Q����VY9/6uA��y�ev2$�?�La����(����UH�]�(�* Ćn[ ��c��*�<�ՑW"���8~-�
��&ʇ�6F0ҊI2ZdPX%&w�]rP�_�qň.���0r�YTU����\���F��?t�T�}��'�!� C�\:�2����4�%�4���U�2�W��`��Ld�i��H/���tkn�4,�x!�Y�I'�O��^b߹6�M�ēf�� Ӈ"����~,XĜ���V-UJ׈��β�v.$�<��LTLaV��UiT��J�'gi��N���
�T�w�'��It�4�UV�pX�݊��j)��݆�1��ы0l�Ц���N�,�a�v;(s�b��-�i�H3yy+�Z�E*�~���!�m�1�ɖ�f�O��L�,��Տ��)��R�&�z�2�*^a@�>AWe���byn�1�|s�eT�#jz$�� ��B��_��?h�A �X�-��ST� � �����nwO���n'�;���*�F3NP�sC��E�77 r;1��dIcN>ɓ�l���tT�)Z�vh=܉�����Ld��mH��Sub�TO*"|0J��U��+6߉?,c�-�,#G�v�-(�9 +U�fY8�r�ћ� ��5%���:���|M<l�jM���^�U&̯��aN'�Z$QE���Av��X�u�M�*�4U'}�}��1���-��@k�u�;Vb��I(w؎�RI��>0�i4H����Pl�ZD4��jsm���ܱBj��kW�ދ��ƈ�9�X�P�Ϙ��CoBy^�����;����ș+��̸�zcRAZ����7v�1;��EUkY�0����ѝ��q���lo1O� zc;�ɼ��%P�g�7@����+BwV� U��K-�P�W,��B�aMS`��B�}*�y�r����h捴ѹ:�O���Ԇt+ ���e��1�,����;�Y�B
(P��!����!���r`�1��P��\��mQ�F.@h�E�K}e,����+�%�-�%h�s�^i�,����`�U��  b�"��W�#�(���ī3F�2��[����c��bx�H��$<#�(�_�	B�ĝ���r�X�ZI jr����+�Y��i����7�P>�O�Ϸ�¡FC�4�pzc��#?�YN+]�e
v� �=1����>��F�ڬ��$P���'�w(�c$tZ��Q:P�2Y���b�μ�_��o��O��6$���oܘ�AE��D���4g5U�� ��
$�)c)�;Ԛ�W��%Tq��FM�oڻ-Q� r�}1�)'����u����] <�fU<�Ke.�w���<����6���a�f�G4Wv���v<�`=1�,)d��1�cĈ6Eb\����3`�m�,`J�����|!�Okފ+@��?%�����c��0l��V��I�t"��J��P��v���Q�c�vM���1�DX�G*Π�(�,��*�P>,Թ����#)\  �a��xՍ9�h��&%T��2� Rl"�X3t�d�De)��G-���s�E �)P��~!B����;y���k���S")S��ü�ŃF�UB�Km�U��}[�����ɧ���4�/ͳ1�PW�i��_(	�e�@��R���),g#{����|qrخ�-Be1g�4��S��o�o:3d}�G���ːc9m���^t�q�ζ|�\y�I�cC��LB=l��vR�s��3O@��ԡ������7�cÎ��9)�c��u�=>�������W���{�ѱp4.��WP~�M��E���eX�$2�)��Bh6V�� .��=�N�:m�5�.�X�Z�z�ģ�K/#P=v�\/��~��틩ju�t'�������[sir���s�s��??��Wi'�<��Wt}��$/\�%f�s4��@�Eė�b�#�gż��hOۉP+#�x�c2��Y���������[��v��Vݱ��WP��\r� �Ib8�#����n��ֿҹzwRw;�#��/��f��tV�$��W%��WM!j�y�b%�c����z��};0m�2^y��WJJA�y��ԊA!��!��\�^��&�:���wN��u�sjs+zG1!n@!���x�H��tvfV�uƅ��Z��V�Z0j��S��ɉ`UK7�������t7m_�..'�xv��YY��O��� ؖ���ՙ�� ��K�C6+ɪ.V!K-'-.�	Zg�!La�28�4������f�7��˫��?����,nP����ݲ2�z\̨8�/Ƞt[����Vc3�Otl�bNϤ�!l��ȼ��#��&V<�i朂#- f�]K)f32�oE�u,e,�6�*���0�!Wl�S;i��� EV����ӝ'��8��L��L|�KFk��7L���T	���rL�Я�`� c3���*)/�-
�Q	��$�K�Z+ �Q(�_/���P3,h� ��$%�
�_&49���+~�t���L�É��92�fW��h-ҁ�i�AS���U>j�rQ�����~)��P�{�-%k��Dd�����@�fh#n�r�B@NL囓�1��Z^A��f*ZloG�K�/�	"�Ê�c�Q���_�1��
�`��[v��dZd���ڟ]�lT��c%GMa*-(��lqR�pT0�b����� � ~�r~|U�R��"��*Y$�mvP՟�ܐ|�fb�M8�d|��v3f[�A�/�n� �~�m����$��J_zE��ܞ����� �!y�A^#��SXȱz�C82zE��]d��h��'�]����"����� W�VV�=j&��^SF'by3C0UUc���K�wjA�&�$���@i����#�7�oLc�N*oi~E� ����2hj1㉐>gGr�r���vn,�I���<�d�iE��~vNd�:��C[��K�A�zc��<ً��k��f�f ~�#�o��a�Lc �|~�Fj1�9?$r��.���VT3��G�1��H��xRD�L�AK�`X�(.Y���?%�9��':I�̇u�"�Z�ǣ�㺸�Ay� ��w��
�3��f�@�n�,��M7Z9�<���n'�<�%�������<���ej��x5�l�����FŹ���Sb��nfw-d�?�`��VÀ�l�N��a#�� �Ȩnu���f�������ոp�vtngLcQ��cq�W�
X�I� �V );8P9�ŉ<����QJ�1����P�	L�mǑ|��.ʇq��D��V�6,��BI1!��h�k��2��V.��ZTQ<r��]ު��;)b�o�bv��clE��FJ>2�]a4,.� ����;���c�b�3�Qjo�Ū���Z�]Ԉ�7�Wk�([Į�6�ZA*�*�|���_��>�y��s_�!IP%߾6h�E����>;E�+��g2�y�C~6B��m#��hQݹ�^�"@��._m��Cog�]k�9��=����ZH�S����S���?�V"�@1X��Y���N��a�V�A�Ͽ��Sr�����Ft�?U0�׿�	�(#�IP@!_ȍ���g�����!�U(�)K3喊��Y����x��1o�Q ������}&5�R�&�8GJ�Z6#���sk��R�ٳ���k��6��S��H޽N�=)��3k�e�F�}�
������P��p��6��D�.pK���B�����X��/yJf����l{*�3؆>��NN����T��%�p9ic��&�w(���7]�౑�-E�;�02x`���cgxB0$Z�dZZh�~A�N�S2.� ;o����f|�C]�,E%+y*F�F�#�S����6�-�hqj�/cʕ<&����� S{aZ9oa2$�ڍ����c�ȴ�� 鋬�@�Bc�yq������&�Bc���ӓ����OZI��-���z��$��\+���;D�������"���}�: �Q�"���-�?(B����U�j	�|��+��'Y���{s{�d�U�r��无�*��|{�6�E^��p�+f��bmā�p�}�f�k��=R�ؔ�����u�:R�z�ʗ��}��&?d�T;b�v�Zl04�<%c0,�����7?|�/�>{+�d-����* ��%��%�Q�"�v�B���씈�`K���P
����s�e��V�gy~'�3���4꽐}a��ٰ
o��{AH1�h�|Ô>�OFK�T�'NM��C��p2���gv����Q��AF�^�N>d(����+�N��'�`������ZZ����.z��ה7T%�/�:����������1�}	;�*.�9,�p�flÍ,�y$ƣ;8���M�3��}k��<� 5�_��9f��Fi�{]/5�'�e�P]�Ź!�T?zR�A=#�T(���#��/
:tbL#s̰��ȍ���]��6{jnV����Gg@�/��Xz�]{�)sO`�hFaƨ��t�ٜ�Q~�\`�Yt�$�c2WR�����Zu���vքD~-3��S�8li�u�o���!���ȉSދ���v���~V�bTK����~��t�1D��	����B�� CYv��O�����Ǘ�d� 7N��������������b�_��K���E޺�Y��8$kI>˚�_7o��Z��H�����}۫'n�I�GƚA��XR��Ľܚ�(瑏e�b�[���r����*;��qC�/�2Q{�^ˠ���hʼ
Ks6!��n'}ph�M��d����"d�Vjg���Brh�y����QN�Γr���Y�n��mvb�~5rm鿲u���+X%4��Q�{�,�L3���U��m��É]%��l�s���<t����YE$ޖ�'�����]i�������!�d�Ѽ���)�AՏ!M�,.��(�ę]aV����ޝvz�0c�uh�~���sOj�w���+�5�-��T��	�]`2��pCY5L�i���)�J� �=e���7���#�m*������O�Л°�a��;n/��Cܥ��u��H��	�=GO1շ��=5���*��0�[f�Vq+�[������у�c�(XSa���r��=Zb�f�x�)g�K�$���^����n�Xen�y0��.՛rmq���	,D�YqV��(�  d��tB������w^������U=�9n��dҲ�S��S�m���V���|Cm0	�C��҂�����KL�^����k���(��g�4�_�� ��
?����n-��!�
��қ� I��}T�@�3p6�Q�+�l��P�޳�v��q��TZø���.�U ݌W��k_LB�{����줟�ՅK9w�o��W��n�|{��H�SY�JZ�}�T���H��z��/�@�^`�dQ��6��\��3##%Lt���R O	�G�ž q�i�����
�G6�)ٱ`�5�=���ܓ�q`8m�1����]�6�z�r���@�d���wW<G���'�Ztl�j�r3̈\��	&C��]�(Z��HLrdL����RP+mܰ�rY�ؖ�*����Й�*���C�I1��)Rv�y�Q�LP�N�B3K���}�[������)���æ���Z�qu#iC����J�&L�����OO����_s����Cg���9XȽ�'��a2�(��Q����2"7�^S�ub��+^�����Q38H��d��T>��;kq����� ��M3��7V3mly�:���9kh%�`(f:wp.� ;�h�_�F+a�7�VP~6�2s�ӕ��Ѹ)~�ݸ�Ю�X��XuQ]��֎,��t�!�.���)f���6@.��s,�q	gLe��3�?��a�kl��W�='�כ�24�Z�d�7w�_�2y�_^~*�Pɇ>q�m2Q7�,.��;���W�Z �����.�[#\%�I�fO��(G��SvK���Q�/�d���!L�r��"̭�5j�����2-��:$�&pNdT��
��_�v@U󚓈%�~����{�OM2��*���? W�0H�.��bV.VO�@��(F�f��/��]6<���;�Yz�h�x_:p1��]�*��&�w��I�?F��~x]I���G��	+	�7��Y�R+?C?|a_��N1���C�0��?=�������Z�N��j�ȳx�e�׿og�Wha�wr�f�t�C=����f��GJ֡�7=݈0O@��D�5�K�,ȷ�|�ƈla�bD��?�w<�׶�)LV����$���r.�S���[�,&���?@��7�0>�|�I�b����p��'�Ϸ��ii/��љEH��"��I�y��$@��)l��AY\vP1y�7��P��CA=	}B$G*���sK���zai+�(�r��x&!M��z��:��#��=�*�p��v]e?9_J{R�n�Y���})�*��X��w�kL�^ˢ�]y�Q{�c�ϊ������WL�t�9��5�vM��Z���d�<k�;o�W��������us�l�4xɖwJ�H����B��)[�{��Aݎ�7�Cr�����}�r�W��/�M��:����.B��_x���}| *���B��9tE-M�V��<�8�$���|f�b�l����k4����h��͉��n��R��,�Ѩg͝��r=_\S�����% �O�i�����=��s�*UO𞩣ac���0��;�A��L�PW1�����q�Q��#��rN! "f!1^�'p�Є|f�|�k�vNEX�Z����v>���Mq[8{��h��wq�1�Ë�����Yi�-�Y9�-䀙�:��,:9.����0�F���Um6}�_�-Pb��HB�X��J��WtM���aK[�8���0��]ϣ}�ZPX,E{:���5Y@�U꿞v�ɳ�K�ݓ��,�e�a�����F`�r؎c�\��F���t��,�ׅOc�9�˓�h/� ����I����*�֚��~i�U�	M"���_q���#EvG�t�d�����r��Ǻnt����Qhщ��8XU>X5q�33���>$�{[p���P����p�U�*���	\0����B0(.l����4�*�^��Zҫٍ��9�&��X�#���/��r{�c>{f��r������~K�n��<�򘙤�z�D�J�eE[ѝ�9w۲���{��$��!�b9
�u��X�>�.��H�<�_6̤h�ߦt�ȭ V*[ޝ��T�~P��.5e�Qy�r؆I{��]H����; ߙ�ݕ�G
�K_E!�_�ڲt`�a]w���KjT��Tn����v�����8�7B8k�o�\=E������V�"�V)B����;@dH.!z�z�b-pJff��mUs���������o��斢���&�Z8�M3�Zk{�[w��%�D�R7�M��;v�4[WPr��,���fN��BL���#�On�N(�6��1f3���`��KZ1����r\����ؿ8E��j,
�b>�8��;T\}������O"ŵ�k�i��w=5�/��
�
�.�5$+��ѣx�VǱ:�kk�Hꮥ�YIxe�tk��o��Q�m�~�u�;����,�'oW����/�U@u5ģG�Q��H#��2��������_��a�!�b���ܯ(Y��p����� Bi)'��r_H|E�;���Q���8�����;Y�ְ��ָҤ��4�Z�����8/.�R�����o&���hd�������J�o����T_�L�e~���|E�q��Art�T�#'��$f��fg��WC�+dO�O�&�Ds̪�p���S��-�z?u85<4Tj"R ��R���:���	����#��W<@�Fz������~юkT��<|�4���U��/D��U��돪m�)��B^��4�-��̄�w�����t����C�!�d���X��i���>(4fuK��`W	7�_��j����o�.P��� ���+��Mp��c�>�U�X��5Q�!���w���c\-1�l�g�'_<��Z񺧪��MR��C>��/)�r�3(d�ң/���/?�i<��0�n#˻S��8���H��U^��r�ù�щ)CA���u�`���8 ����*�V?��,�s�Ua�xR.����p-�R�-s�g��N&�K�tʼ�`
�Є����2 ߵ`�f���V�J�8p��Z����&�O��������A\��>S�j{�CZ�s�x�w�Q������6z���/1��o��UJ����|��q������G���D����K�.����2K��A����R�����S�3K.E7�7�`CGn4q]�1�\�a��7��..��_T�$|�%��2n���5o������ҟs:>�ЃFN����TW����sѐZ���V�ʧ�Y��
W�Xq�R�&$��@�Kܴ�[qo�)L}1e�'��.��Rx�υS���Vv�c��*�`P�/�D�ɩ��hc���Q�d��֕�Z�gg�zX�~Z��q'�o���4����Lq��V_��a�>(ϻ��\�J��8Ie���GS�>z�#��
j'Ë-�_@�
�wzR�μ�PE��ME���:�tf#��2ɦ���P�VY��P��p�l���'��e����t��_G�xÍ�އNۀ^HR���s���k���|��,�Ք��(Qd���i[���_X�xR�����uzF�����X�Xͩ!������$\��G�* ��[q��#{�k�4���_���@�u�vA��Wo�{�&�N1c�F1���84�p�9JH�s����T��׶�Y�}�)���	���dC���Y���W�;%���Rң䜼�!�o6ߔU/��}����sN쌸̸�H��`�8e�҄õ.�K�V��J�eϻ^k�㪊D�L2-�M�0���X��d�㕯�<�Z�g���,��l߆�/��R�E��4�83v+l�NPp��6��"�6ò���0	�/����H��<>����E\����d ��dZ�)ũ?�����O��]�����5W}(y�cUt�"T>���5,������ѵ溥È"�6z��E���k&e���4��QA�Q��l*��2lX�Z	2�T����z���1%��Y(�����0�Hrf�̓�:���>��������_&>m�)��\�5}���Ȩ�f��O������t��o���L�,o1��Ŏ
�B���o}@Y*����\���D�'.T3�ľU��PZ�%Yq�lw�+��?dP�Fyy�1����s9*���(�/���`�ڵ�6��2-�@�XZW> p��[����0��f�?q�)^X�������&	\�K�Z��������䚉y6�aXH��U�t�K�wp��;n��DC��]a�(�s����D`� �V�kA<%78�}�a�n��A�i^X8���T*�X\���6�cg�S��@I�?����z'�A���"%r�_����>'��(���ނh�5�\+ }�_G���-��J�h�F']e<�HK�\y�=�z��|��2l��T;�:G	#sg���FN⒂�n�·��;6��M��3՛"Y�p!������X�"5����4�%���,���~B9Ck�o���z�I����[&`a-@���Wd�m��'	�����m�����3�� �I�Q\�V��7ujWЌ���G��]m�tr�Oᗌ�	�L]m��?�-��-ˢ��v���;G����ݲ�$ٲ�1=!�M�N�f��J� (��7�3Uzޖ@+��
��Y�������x�R��_�7�Ѫ{�nz��_j:�}L����խ�t2Uf��tM-/ޗ��"z��Om��m�\���1���_�1rC R;���c�V>�V�X�ڃGܜW�_�%�QI?�(��v�+��EQ��<�3R\'V#�~`{/�[4�[:��`۪�o�G槺�!a_�Xm��+��rQ��	���"	�ñ������g_�c�u^�u�	�����,W4T��V��Og[?6����)�C|�vw��t��J�}��q'�(_�`U������Ν$SZ�<$K�<V(��ڵe��,!US��1��v�W�o�Ko��ՎD������\�{�R��#��	t�Cr���-gNA���*���Yu�e���_��K[�&�]�0�"L8m	���rI�H���:�P���D�y�5�D���������j�A��YrI��n��RT�1�2�,h|jSw���`���u�Ƞȩ%�w��������o)����k��,-8�Ɍ�_{y����ɒ}S�S��w�>��sa�A3<��TL�BQ$�+K��I�v����J��\�ԕ�r�:��u�T�=���	��?�=Tj��p�gڦ<��7v��D�IF�\.��E<q�:�Zj\��7ʋ�Q}�+�JoP���rL�_̼�
A=O�V��������Ó�_BR=�,'���y�]�����A�1�E��)��%A�6geL8��A4��QW�L��f�����*��n�_�݁x����b��od���N=#�%�j�3�;�˼��,��09�)Frb幺<�&[�{!!m��������t���X�� �csd����T+,�M\�zdf�H]�58� ����?�ZJs��b/1���}��,�P�:P`��)�N�׾�|����xa����85<ϭ}���g��њnͫ�la��^��ݿ���ht�EOK��%����&9~�LWsR����o��]r&I�@��4����Ϧn��J�챑�����`��!h�&�'�`y��lN�I��Hi�O��/�qrW@ϖ� i�n� �t��GC���C���"H�gד}�zN�˨��W !�V�8�� �U#�	^k�a$nT
U6w�(�ѐv���#�,�	��Ⱥ�7��
�JI|X3;��D!y�5����*�eՏ
��Fv�ԟPچ1�Q��d�뮄�5��z�=�p��e#��2'�}��,�s�X��\�1���V�ďG�~�>���J�wq��U&�M�h5fQ7l�4uP~\�E7I�n?M��0(����T�����O�~|YͤM��\b��/��� V�4V%O5���2Q�:<z	�)`�<	��O,>�|��~'8mLͲ��{�
N�L�M�G�z��!N�O^aٷ��yJ:v�����"�*T����{�9��1�t���3*�[अBc�T�Ǌ��K4��v��O�a�� �p���ȯF�!��-��v݀�7�����|��(��>��������O��xi�F6�㧪 n�I;L�)�1Y5�WP�[�?c�� ��.RI8��W;s�æ�;rz�)����7bw, W�(�V}�K�=s�|� �"��L�2�+
�u�t���0�y�ν(2�9v�M�#���n��/��h��t� iʧ�����U�|`U���c�(����{�=/O{nސ悠V�2��4D�4k����:�F?����s6擘#B��?���kU��%�a[�&"��n4��dZT�<�i��gB����S���H+ғJ��T���W$%�Hܦ/�4
�K�h�֫+�`T0�s�"�,�)�?�{#(ƙ9{��?�)oզ�,M���4W�e~���Hs(�U�.��7�u�S��Ho�z���g����������9�U�(�M���Gt�[h�S-�"3YD�{�b�,��޲���h6�4'}��+r0�H��ͬ U+�Y�*�<���|:��_7����F�1$��t�L�$�����\,�&�Wq�3d��H{��>Τj2�(���m�m^
-��V�N����Ç�:�)��n��N�#��'�K��/Zx;~�2I�yWA�ҤP��[�-��z��w�o��]�7p<���o�"�j�@����Y���<F����LXh[�0�x˛�|��� 2��ȌܙEB����q�ˈ�zʵ��!h~�6)O�
N�}h1�"����S�����o�������VS���V˺�
��f8]3�]Je
6��ſ���1cpr���ns��M�U�j|�d=K�+�ʦo��<1�>5g�/�� T�m�aL9�l��ꭜ7dy�*��h:���EI�26h�Z���"	�bm]]$Օ��ߊ1�4��<�� ��!T��X���U���G�{���S�cu6��� 	�۶��R:�7F=Rԓ�x��K�m��7�!tm�uJ�%ڦ��?&7;H�eS{��Y/��R�Y���͐�F��'�a#��TP�!L�ݗm�X�D���zÙ�5�bq��;�<��x�9	��(t�����J��4Fy@;F���O�ȑ�4����=�/o��df��FX�H|E>��r|�A��of�Q��a�lc���;G�`%Tf�=ۿL ��"�n�0��.�yGW�5����̷�ۋ=�Y�4#�vV�${d��|g�'����a<i���o<�i�.K�bş�VC�Ʃ,��<VI�h��U�Ô�#oݩr�N��RؐXq\�����krz�)���=GL�Έv���|Lal]��l�/�F2�<���u��v�Л�7E+�B���>M�n9(��X�`,+g����Y=]!Q��I5L�XGD��q��J^��6�,r�G��@�N{��t���"��84	iR&3���f���䣏���8�Xeg3a��5	-�T�-8r�~���8qR�B��*V?'{��Y����Xo7��K�CI�V�_]6�.2wZ�նu�����xQ��A���rڲ<Jl�8n�
q��8w.��K��0���N�Ȗ�s3;^�M�l��T�G����p�mZ��t���P-�����o��Q�����`�͜��D�a(5��0����cѲ	�R�KMo���I���dd���\O�4~��)Թ��F�Kˁ����~Δ�x�]y�L��wM0y��=����OO��=���_����	>�9ڍ�CI?�_��]Ė�	$�'���դc1<���F�;JZ
2.��d�
��LG�Ê#nnp����}�����skP����[1����&@��SQ���D��\LlB�	$(1m9`4HO��ډ&T�Kp��[M���r:���[���y��p?]��Z��yJ��}��GT��͛ܐ���Y#8�H��_�~ړ����u
ChvSV���_Q����S���=��A��
g�~�S:$=��T��پx���B�=a#">+iLe��<�U��`��U!�P���c�2>�<G��z5�.&�.�ҘZ�g���C��݅�2u3�h��Q�JǾ�A����@�(��4Nu���f�xB`����y
�o,���m��xsf���hN�������ǭ�
3�ݫ�4K�Df0����D���w���ˇ�2�P�5B^���q��5�kX�T3F��d��������s��b~��uº�	!��r{�Q��}Q>������)^�t%5��I,:�����I�yۈ8��帔� �U���c�}���I1�+;��*87��=KN�W������R	v�e��Xq;\�]3�N���<�<�.'��OE����(���пxض��"�I�l?vCp�8����V�Xb����+)}���8B�!��)$ncv�I��@H�G�ŏ|*�9�_YU>�QXP�!L�4n�$��'v��y�ۗx�×���!��'B(c� ��5���xL��`4M���>B����Ä&���S-����3��|Rz���P�ρ0�P�G�1���7��[�7~(�p� 1r
��{�	
3����F����-���p_���/�BI�6'ȧw:��
�E1�(�>���'�Z�ضV��4�ձƊ��Q��?C�4�>�g+���mV�Nn���.ǂ��ޤYl��S��ɱ��2B+��,a���f�npJ�#���"���Q�^ts�����^�#xW`�wX���Bk,�N�	�޽��c#3�ō�)�?=��nG�<Qh�x�=��;)�e�P�d!&�.�8�3���S,��Y�� b�-0���[���Q��/�)<�Y���E�=��.H����S�rYjũ��G�5�7}�'j�Dt�8Ѭ�^�h��i�u����sǆ^�xTԇ�l���#7��%=�a���f�����p�u���I���J���<����c���^m׋ƩU���EG_�û翾\^�ⰾTl��`z����{3�2y�X��Wb�=�ϿA<�|�ؑ@�Ŗ�Y������(���͠(V�On_P��K�lmß2�q4�߫a�ŋ^��`��r]U�w����XC��*R��,�.���I~��w��?�e��W�LXv�W���и�y�f#ţx�����sp*�Qt���/s��}	���)Z�V�T�U��DB�*;S&i�56סg�����In�V."�cl��C�]��~>f/!5�-��+��u�����4\��o��ȅ�@o]ͻyz���T��R��^����{�
�!n���osB�(��	��Q
ţ0�p��!H��YW�ff�D�G�w⅙�-_ό����(vՏ␲:^�����so>�n@��K��5&S�.g]�sgK��W���~��.*i�J8���1bV�����g(�!�~F��ɷ�<z\q��x�c��B�5c���O���0�{�է�J��}�(6�G6{�.?�/s�;����Eaj�Dwc�Ɖ���e���O�8�����\��I�u%��ݶa(��E�{e?m(s�i�D9 �owr�/5&��1߱Bo�g�C���d9���] FE�=��G+�rQlxʻ��auc�򃾕v?� xgnoZ�q�{�:��[煩��d#D�>��d��V�M��n�a'hP���� ����f1� �	@Yv?R#����E�Ji���пȘbds�V=E�8�ħZ�Sk�o�����$�Ф�R{2��]�F���'��k����r5��$c��*�v:��M�r-ţ�Dd�΄E1��� ?{�)zD���$r˥��ٺ��5Y�j��:x=~c������#�{���i�3�-1�������~5�{�z���^�p<Ʈ��`�{/3�:��*�
<p@ױ��J�.�{��n�\9��sH�o�7V�*2	��΁�ͷ&${���<�H��a\�l����]yΉ)Ni�@|�9[��m��%��d~�f���r�O�Ę��f��Ŭb-�����,����Cq�؈�+R��}'���2z�W�
x�yy5#>�A�馨^�j��z�ʺb���I6�jm�_���`C4�(�&�����<�3��;�<K�
]�j|���D6�=�����o����Է�3�)��߈�峸�ȇ����'9\���z,��?U�'ɝ�c��6��?/��N3��0^��y����i�k�8�BY����s�D,�\kg��rjc���5���:�4�5ط�S9���u�q�ˍ�S�L����B��2?C��s׋=��F��M�]�F�W$TW��2�\�1���ˎ^!��0��8S��+F�/}Q�i^�$d���v�R�Y|b[%8j�Ë�Y�E�����Q�F^�Z�&����0��etWJ��� ��_�YQ��,`!�Cqpwu�hp��8�֢��8q(�k N�>������O��{��� ��o�+�gx�6�k}^ky��r����o�Ovx��,��,@=��\h�Ș܀=�3K�,TC�V��}˒NIi�j,���[Q8�WK�Sq�:����mo�fe2|�L���������je��*;��k�
<�X�#Dɬ���.�Ƀ+���/�"���ح<���f����kkz�a�a|E�1πl���U��ש������&g��!�u���%db$�E/J����c�Qɛ�*��M�Y>�]�)����w|��ׯ���={�_�*^C��Εߡ{� ��͏�fs-��BR����
���v/Ǿ�m
��m.(^;C�[ϖP8�Mf�HaP����RG4�u�eZOL[�MJ�̗�r|c5������N���I
R\��%N�Mz�b�������ɇdm ��8b]-��9�(�yJ�tVӕ̵':���I�wN��I�Ԏ[e
�=�L����'B��-��s�M��|�@Q�~scy����@TV��a?���"|{=��Nf&��T���
xA��oS�A(Z'!h��b��N����'[f�R����t��,�ǰ��~�Ϻ��v���i92�.y�daS�$h{z���jNl]��\b�n�j:db��V��ė�<��u��4��ο.�+�Lg{��6��f	��^#�TWWҰu�=G��F%�������,EI��K��Ҧ��X;3"��+t,���*��Ȇ�XE7Hӏ���X���77�9B�M�{���/�$m��b����x���Q���B��p=������g7���xyJ&���.�Ã]�Oi���
�}�q��j���d�vL�G��uU��3^���2"�:/�\{\�y#8.$��0˵`�z4���O�Fz�r���BA�v/��~����S�sz��4S�U�������Pb�po�u���Z����R�] ��=�]:e�뿊9�O�����iw�{ܥ��l��7]�-)����"n�y���u@,t��e�X����ǎ�Lȕ'I0�g�z�n���bZ\ �K���@���&��0/���S��ԐB��3�?X4����A��d�;ُ��c���_�Rw���������V��EG��{�Β�]hyn݌(]�O�^��(�B�Mw ;�$+(T*\h��ʻ���L˅��J����'*f�\�YhA"���+̛2�λ���n���y�͕��b���0�����l(�T.}��>�=߷�E� �n�/���Sm̼f7a�2�B;�K�m)-�V+}	��,�!
56�"j)!�Ԑ4;�g�,��:�|o�E����d~���3s�h��M����弤Z�|d���\j5>�6OٸH\r��	���]mD-��/���[�ҫ-��߀yX��l�G�C��a\�c�U5eݮУ�����?<�#S��i;�+����!R�6|=��s"1郀 �T�T<���t�����F�w%Mx3 �x��N����g����sh'�=ko���L�f��WW}��5xsY�s�e����P�� �1��w!�`,C]������hΕgͦ�l��}�R�s�|�`�g��hj��h�-UjH+n�+�9p��7��=������ܴ��4��	�3�a��c��\�A�{�'Z�.���{����l%ѱ�|���������Eùԫj���0����82@s����@�pR�UX�jU|���d��)�&E��5�����TG����T��L-gg"�wr̰�� d��v�Z���p�|��	Z�Sb�tޱ��8�.�Q8����Ĺ@�Y��]�ix��N�>��ٌQ�����<�L�	��0��!Irx�^.� �sm�=1-]���7?gJh��l�r�Ŏj�!�v��яT��X�7r�,�t�v��S�F:�p�0h���HMnۛ��I�Jvw�>Ԝ�d|3W8�!'�]oyق�nG-z�D'�cZ�,�L1��	_��f��J[�.��Y��X�SӃl�?�VVM���(�vѴ��8A��wj�n*���;�G3��}���(�R��*�#���a�زQ;)��:����U��v��0a����T�Z�$^3Jl�x����M�<��i��|�g�pH\]{�2@I�P��+�w�:��H�mk��>��k�1"�y2������L,�W7n�ke/r;��;�m!�����`���g����]���Q������0~�JuC�+��6��\����L���a&���N��c����#�=�{�����kLC����,:j��Bh1�|O��E����7����K�������<�,0�Ŧ���yp��K�������#ծ�a)1����j(�p�L�,5�x��T�ʵ0D0Gҫ~z�]=u�a���])�M�'��Ţ�ǔ���.�f\X2��_�Āsj>XD�J7�y�B����3���Ͳ�om�>�x8EZ7b`�kj��R�2�U����z��'-�4�|�\M��zÝ 5�Aw����g"y��{p+n��η��o:y/��&�H���ʁ�=� ��4JO��y�7y�̺�n{`D�����r����o��SBL�8ì�wXKh��8��3�m�]��k�[�����.2���x"3�G�1tۿ�q�U?*z�U7���XsD�
�f1���&��䤡Aw �� �t(%���4�q���pA�順�� Ν?pn����}�9��{��Ლ �d����KM�s�u� �|�/���:�-Ft������.�q��F�at�I�M=f3��e���%�� 1���	c��iv:�{�>*��?M�̛��U���%�9�!��78���f�,(������%#.����v�����<'J�E�>Br��A���$��n��ڏ?���$�<��X�<�1�O��G�C�+�,�J
��D��0ܵML��rΛ-��џgC�w����P#3U�9����C��=�M���٢���D�����R����"�j6����K&Y��Nb�ͤ$=��:
O�c�n��� �+~d�U��&�mT3�A ��j	�{�J�?No��(�p�5���J��E�F�XL�X�Pߊ���y����drּ_A��VӢo��;_v�8O�'�J�ß3X󃀬���+[[�T�?����f�+� ˲tov/� ���o�c]�xr�Ȕ�]������D*���$:s�u��@�`-}I"�E��'p����=�s"/���M	�����:8���L�cN��!�aE�nB�q1s�h���WR�kXg��.׫|~���`����5&���>�2&x|V�h��S���ą.�7�rb�S����}�F<�L���jYr�'쵪�/7���)���*�LXzRd�HDAi�P��p�j�=��(���a�*Ġ K��f�~97�j�����#�i
:��p֟�
������c��N�X|��? ���2X/�>N=�h���J
��gFg�dn�o�^ ��\��I�j���Be�0%�	�Qɉ�%�=�J�[�����Ge���:�mc�G��y"�c�S���(���ȑ��-δ��[u���Uv���_!��PY�&�j�_!|�6O��Y�FJ���zO��6|Bl�~��_��\[�Kp�=E�"�)`��ĒZu]~�o]:LФj'��2�v�F���#l����eX����
�����	�T�T��b�p�ٜ��w��ˣ�bUP�����j	1q|�u��k"�Bpc�V:��9e:h�|5~[���@wJ���3?N�"ۓiF�-���EG��n�* .����yӅ��-^��h���?l�)�y	�.��ڋhJ�����=?���<vH�����麍��b��2չ�Pg3���W�̇s�FI�������pk�CF��=�C��植Tq�`f@���HR��8�4kx���b�F��"��j�6���A�\�)�A�4dG��roc�6� GC���v��@���)����I��{�N;�ی�d����˲����i"3��(��"��ϧ�{ԉ1�k�����\���_��4ǒwox�Q&9�i�=<��`4��c��,���0�����g��x����{��F��{��%1J�l�1j�Ĭ�k��j�E�n���&-*�0�O������Jr�=��~��snp�
ۧ����
}������@�$��AU˛�M-��)�u}�I�$
�hkc1~I����y��z'}�MYqW� x~������[��׻}��qQ�?���+����g'�pau=�A�C��û\$�I�$��su=>Ч ��o��LuT�2M��ƥ�����ԅ�d��\���(Vލ`�ȥ�}�b�ac.�2S��V
ѫ�1w�4�Z�����%hV&���o5�쥥����Xv%�Z�X(w�N%I&:�5��A��Za�\�8�*~%�_$^6Ձ����l�e5�c�(�+]O��>=�����Xb� ��љV/�2�=���$Ў��p~�� �%��(�_���rG|��)�;�ҠI����lwЧd8ܒ%��>��M�~����a�2׎��<P���W;jR�k�����}�K��Ǒ��D.���B?8�穿m��Rp�NM�UW�[�!��8��+9���T�w�G�2M����O��AGbq7!�'�L�+�8��o|76�ZlC\�7���_��7�jD-0R�f�B>C޸��L�b�A� ��}�â<E�R_��ۨ��5�{N�[�G��w�F��j,�{F�r檼��k8��/�t����w�:!de� {=y��|�����N��d�_��O�=v�O2�ǢE�gQ�nX�[�/Hi^�}�J�Ԏͺ�&���Yl��>����!?�_�qi�~��YU�2�6���.e:�lۣ.�S��T����9����!��5:�]��/-f�્?#���4���y�R�/�`d�q�/==LY}�_mⓜ�խ�!�A��5�cN���P�N���gW���᠕�e.Vq��D�� fZ���a}��m����4q���R���y����o��]_�����qΡzHB��e~sxR?�u��̴E�ߥEA4aߎ���l�����cP�D2u�T��?��H6U�����Ln���4H����w�K�����T�<�������9�Qw�f$<wO��'\y i�o��I"� 9����g/0U��TF&G$���-˪��S^Id��A�];��y�
�S	�< �D:���$l���uRݏ��n�ϛ���B�S�je�"�]k�[��Wz�rlk5���>�K����7%�j.J��-Z�~�w�z�
��A�K��{�e}Ov���@pG��Yܥ胫x�[�t�zZ�U���Չ�S�a���ϵ���}hR� خ��F��"A_?����V�`�����61&%i��Ѥv#r���n��(ix�*Î�"ߖT[}U3�N0� $�G���/���1�1�(�Y��ˎ�!;�?�J��0��O�h\��ú�j��p��D��)�y��-IY��5^3i�+S	�H���]��	��!0��	�){ԣ�jH�Ƕq0,vN]=6�� �_����@���W��4;0{l~��9S,#�ҮeRЅ-��ب6;�>�Q7357�pN���=��!e/3��V}`����UvfweO����W���_g�u���}���%4N�0�8�|t�Ǜ9��q���T��[�3�U�d؞:s7����Zi�,ϮOF�8����`=�|z�B�g3g�uy{��t��W�+���i8YO�1�Bp�{O9Ibx�G�x�B�`a�B��Aգ[4�r�����p]�ܮ��f��QQ�{pY�r�<��5�Nڒݷu��?\S=�� �'>������&�˹Uw�'@��K��^�X1�a�HJ�+�`���a�7U�f����?Y��D�1hcnB0�W^�n�����}G�k���Ϟ5x��r�B�2{��wٳ�w,f(Q���-T�4����ҝ�Эf&�S�Z� �[��p��ۘ	���rv���8i��y��(�p(�S<O���"���qo��;�ZL,��S`.ہ�ƴ:�U��o���D�v��w����3��Ɲ�bt��o�_����:B�K`�<���0��K�6 ���������p'�ѹ��v�x�؉:ͦ���|^�N`��Y� ��C��uv�J5XSv�׵�x�3V��6#�O�+OgSO*μ𿮐3�:�"�YE����<"a���Zf�����U��8��i��Yj�i. ��C���T�� ��H�/W�}#<�!:ޠ��n+����+S�����%�i�;*omw c ����D��X�[HV���&�WS[D�
�Y2h��BC*K�c���/`1��yo�R�����3ىzqO�J��=�9/�v=���G�N�����RB�|D\]71�+z�e�9�}�������8��P_��~��y��Մ�і4�6��K��[j�������i���]ʨ�?�y��߼Uϒ�c���ݸ�OͣPyա��������F0��*c��]��au�>�V�\��a�.�M-
'�äH)��e����������8��ޅt9?t�-�"����S2�$θ�`�XS���'q*(�[��kUF� i�;<%����:i
�YϝVZy�B���@?Ŀ���!�����n�1�CS�='w���I��j��,cLu�8bR�@n�tn{p�����] �ߚ�G��+��=��{쌧���*�9�\w����ƣ^8�g���!p��,Վ�N�����/	fĆ��Ll�|��s�y�%��`�P9������$-��lk<5��亾+���K�f\.�񌚘]E���ި�k�U�C����������|��ֺA�-�t���Bc�@q�S����s3���X��=��:h�,�̫e��s>��P�nu)��/�G��v��<r�K���{�ӫ���U�S��y���!,�q�Q�"g���;�z_T\Us�@��x���!�>�=�K�Gx�*W�ˬ��<�^�q"G�}�\�[��N�1ܺ�Y��i#j�2���L>8{ .�j]�2�9�w�ƀO;��N�ܟ `I�c=:���Ȧ�����k���l���kc&O�z	����I'�?`\���w�+$�X���NTĵW������o�K��>��m�|�m�;�f���dȌ�~����՛T��|�:�}���{�Z\Л �̹��JA,Ey�ʆo��f�׮�V��oi�C0�LR�R3���)��j���*��P������_�[�����*����R��S-%2	io�%�UӢ�U��y����q�J8@p>g�B����H��L©�,�)�,�����T�������~D�k�w����V�|��������OQ\25�>?³��1��5e��ڐ�a��.�UW���<rT'� b�=t�y��6�gB%.!�z�^�-�U)�!�2{�'v+����4��Y3x�g�ͪb��c�Z��%��. ��N#RVFs� �,��Ì\��+Q��{��3HA�͏V�K���[�?���H|u����0���.�*��	4{9�$Q��o$�|����!�i�7����Am�����S,�ҟ`�����S��t{��CCC��v_C�S8�ک!��cE���s\ak������
%�y;D�`���J�,�W��#�oUf%�/����f��s����Rǟ�йX�'�:�.����t ��o[��	D{�ö2�#j>���%Ѐ�!�<�_a5����8F��Ө�3�K�����_�м��5�Y1��#�|I��>���Ś7�)ܧ���r1���pNk) ;k�s(���n�#�
�ST 4�%(��j�$'C&D�D-�Ƥ⊳��ם�h�BGz٣�E�i�P
 8�St��������1�lW�S��w��l�c��}��Z�b��}�Kըq5�f�7����{p�,��o3Bn?% %����������TS�Z�
0;��L���[��U����k�
�6�~6$F�TU��F� m�1~AP/�.3t��~�(�.s\�V(d�sp=�+��|q����{����淜f[*~�&Z=g�vb?z3\9�m����e����|?A�-fpKK���F�*�/S��~I��x�p)�3Щ���=F1����4Su�d�O@y�m�~�4$�ƵL��mO�]��}ʚH�ϐv�|#�:愮�Qj�-�h������gE�l��	g�˛aG��|�Z���Yd��p�v.��t���z�Ƌt�ǝ]���e�T�����&�zԻ�ߋFo'�M��X[�z�(��~f�e�=Uu!��÷'�e`�Ύd�:_}�(�%�8��Ȣ��l<��V�}չ�#޲�d>�y�\}GE��3I�
�g�Y��0қ��z�znL�3I�X�?Y���Pi�a_2N�|0)�L(���WG~���3b!eV<��~_������;Q�#SA±M$(%�~Y�Gp�Gu���,��-�OV/ r��������,�y����P<�Z��"C�2t �^
�M2����5�V[ȯ�rO�Om�XL.��m!jA>��'$�����3�qr��'��Yg+���P��0Y�t6�'����K9������W��o������-���-�)� ��r�,QF#���m{�>aʉj�H��*�Z[?�?99ArX�(�֒"���47���9��+�E_���T[��%+�.�X��k��AiZ���6Ƽ��[bԚJ�g�:�ߣS{��j��)�o��&��ƽ6�%W觌��Z�3�#�=;)[Z�М_�:&��Z� Su֝؟��]F�k����Bdr{_���7�4���dd�M�8M����c �!�kW�L7W+L�"�4Ic�J�ȾW7�RD��1̊�N���p��������dܹ���� ):+-[Z	����	DnVtn�7M��4j-fqR����dL�kyo�ˎ��|^w�w|�e�C?��S�j����͌�wçX��-�x����K�-�d��׼��M���65��h;����S�9�\|Gd����H����Ƅږ���W�ɥf�T<�l���e�go�^2'��}X|���B�2�*�cVd�buc�6�_�����"彩I�6Ŭ�[��w����7�D��_�lf.�
������.�T���/ BA��vj���ג��i�ib��@�a�D9f�D���
J�☼������C�Ճ��\z4�rC$^3>�
�V��wb���zЎO-�M�l�~�t�V��.��$��\^�F��`䁱8"��>z�_GP�����O��
Q��1�?�:�NJ��\�W��g~Ǽ�O] Sa�_
sqY��.�|��UR;^ʗ�h����6%�J�9�ž�N��R��G�̅vFO��/w��T�]����e���Y��b��JP'��^�5Ng)p�E,Z�<W�S��R�t_���OO=�,�����I���ͼk����a���i_6��a*s��+w��-�<�8Xi�?!���(�=ѷw�L��I�0��T��^��e�RrR~��XY�p��t`�ˍj	<8�{wl9O�=*�~?P�ϱ�/ «��	cym�adv+/�_c�UW5��H��c�'�>�BB�2��{)k����@��J�������f4�t�MHҍ`F�>�R卹�������q�h������_�yg7�����k�:U�޴!Hy''΄v����z��⮠�ؗ��O6S�T����"=#�n�����B�U�����J�����I�
�����DL2����i"Us~�p"Q�@q�pMTꇦ��"��͠��C�T�f��o�]f>θ��$	��쓊39/�^���CZ�8Y�9�*���C��P։T���QAI�;���u��u�I�e_w���X��w��[�rt����՝wy��[��'���[	��n�h��Y�Տ?�ړ���pק�u�O��*�ɱ����?����Ƹ]���F��bde3�<ԙ��'��7!�V!ș�4��otʊ|i�y0@6�Ҙ9�?��a�A6�qnЪE)�}�Mm{:�����I��)��2�����}~���D�p_ 
�г���t��ʱ��// Wu���4��ԫtp���̿� �Y�K*0l�w���V��8�	�caZ~��o�]Q�w	IWl��3	���v�DJ��!����C� G��8����HE�?ĚԜx�Yztg�K�gͺ%��ȋ�W�]�K��z�|3u��M����#��@���]ܸ~�����P�k/�"����(U�Z!�$�a��e��ܧk�\��e��ӻ�r�t��o(h� KYy��X�oup��>k.l�'U�$RM���r�ܧdM�s}��3x�i�3��x!�-Ԑu�̖���:L�k?ԏD��u�}�Y��=�����Q kq����i�����5�#=���c����t��-���5�qNvp=����yF�YZ��K��7�^^֘�����t��~�8�4h6�\����.���MN(z�>ScXF��ؒ�qB���FiY�+�����q@qf��"Q��4p=�`�^�׆�PA���G6z�՗rݪ���"�L���-��m�
���G��X4s�`���}˛φu�pH���l^��J^��E��2d᳑���_��L�Y�]�6� ��Fh��
���J�P?�ř:{�l���F��Gi�D�h�I4��݋y=�0A?PR/+�D����O�֦����;�:z���Q���ŤN�7K�Vê����qB�t�b9����S���ˋ�O+4��n��1FAh�{�@��V��v�h�%�����c�\˭�s[Pɐ־�_��>�"vV��(1$E�L��\I�lϔ�i��D�>W���Hsz�0*r·��F�O?�4�_����>9��|U��:Y��ʾc�zf�jƻ�R�0x�#���&M���&+[���!ࡁ.>�(��*"�\�}L]����\����N��E��{Sw�<;��q���x5fĽ��BK޵��m,*�O=B�$`�6\Yy�JdJ�I1n1��$ÿ{����`bt� ��@gbd~�Ģ��~W��A�:ur�6��ܲ,�Ҥ`BϮ�u�4S�	�n��&ry<P�i�Ai�q%)^N�U�Ubi�{��8��r-�D�Xp��e��6���	�L[�����(���j�
�?�)�٤��p�Ia�6�+~p�:�S�q\�w[���@����#c�|]���-���-��������U�3t9#�E�������v����*��7�;�n�m|�h%���]ui���>E�b�;-T���ԛd���Z��)ķ�ߜmFE�x�?����ZP������]�lÁ����[�(���{�+�=6	k�S3�����vd)�p�����ݕ��8o�%� q�p�գEP֤��!V�Ȥ��k|�$T�m�G��"['��M�����6Z��:����j4����w�.{��Ň+�ZS�X�Z�H��?DTy�79V@t;>gp��	t��}SW:��H#ͣ����{�^��S�_�K'&�fm���Z�c�G��V�	E�O��X���nE�E3Tj����t]D�(��У�+y��T;Qę�f���.x)�Ga'���% �3�b��w�����u�*sd=��,-���R�
���S��@]�J���=�1��/�9��gi��r�I����Xx�n�$���T��ks�ʳ3`�}}�KZF�v�B���|߼~d2���~�����
�A������O�^�ؑT9+����9�^�����C�����>G�#��W�ՅR��\&��Q�O�O�c>ي�x�M�߫`�8Y�hd��nq�m�G#�dRl�#�J�؉�u�����ļ��-����Z:�3l{�o��� ��<�^��9|{����k�����ǘ�XFJ\%di�MfOg�%j@��v@��uާ�X4� :�U+�U���MI6�� �>zR���l�{@G�2� ��l�ӢŒxt�ӿ�/֊�q���+�I�ώ�{�$IF���_-�AZ~F���S��_o�e�o�YOݼUKf߹ ����j��8��;�\¹����E��z/�����a�^���ܞ���~���bv�,�`�_ h3�m:ğC�;�<9e�D��וR����^����4z�_)=JT[C�k��L���X^~���Q�_)�﴿����==\��e��7 z���+S�iP������Wk�ͭ�3�ߓ�Q-�ʒ�A
e���؛>�	�ɞm�7S�0V޳�s�
����Z@�����\� clhoQ]�3�f}U�Q����5ip��=�7��)d��BWZ��hj�ӝ��Zl%�Uj�W4�����W��S�UbFE��#��>�9w����u��B�thn$���(�JO��W�X6��,�P�HYi,&*���2Z^�zD��@���s4�j�S��>�݉�D�MH�����MfOڲ���y��;�O�w?��ÅD�b�sb��[���w���ە�GO��o�Pp�)I��=�����}���>�j��q����,J[w�pNg�z�j�5�[����0s��q��̬�s�T;�^���>�`B%�����y�*o�FOO���=~(�CA�Ķ{�®�c�����B�VY9=�dJ_��N�I�\��^ ��j�.��X�� `�a�ʠ�u�Wf�o�?��"S�m(��������RV��PY��'���$���a��R��шv4d9���B�����\1۬����,��3��`�:���?��䬉z�,�r:F2�[����Ε�����vԞ�+~���T�,��18��l��uB�WԵ��-®������Q�7�ݳ��j~n�}ks^�.Ŭ��|�lH6���;�fIv�ԕ'��"�/7%�Ob��*���C�j�e�Pm���>� ���Y�����r_cEN���,��fɼ�.�}P�E)~��$��滹�:�k�ʙ�x�1 �1�R<�����?���s��[��� !k�v��HJd��ۼTQ�Y�8oY�`A
��~V��{ٔ�K��x��wd-Z��;�԰+M
�`�My�A�6��"3%��|����S�S��e��qR�c�b��u;�ѭҬͽ)� ��^YI�W�G�Ǭ:�LȖ�P ��YFf���֍�QR�H��Eީ��P��N�R�DY!h������
Ru�v��L��j`����&O��2j��4*��������]Q^?�Gѝ���oT{Ay~��.i�6���v|Pn��L�,=_�}�TY<L���EAY����a.��/�&88��ʜFUn�3)�͝�_ �G.7ϊ	o�r+�Ie3�H	a$:�o-���}�~R��y�&����喷�+Gć%�  ~�!,-�r5/ M��p������'���c�悀bx��fᐜ+�ٺ���{��M��-�Jn���s�dt�Y��m��&���ZW�^��O@�� �'M,��Gu<����z��.�Ji:��!�Վ�]b�82K*�9弽�� Z����ȺTZ:��$�d���|"V&P���"�M���3^��L<2�sW8b���`xyA�a�A����;�p\ �OO\;h3fb~n���A7enG�8�+,̓�$��i!�r����l'����gr���L9a=� �I���;���x�l����1�� �Q'�v��P��E�F��_�M���5�aӁ�eI]��(��ڂ�)�.`���%�Xܹ�k�=�g�{��[4
o�Xm��#7��D�\5��tp��\�p�Q��]�����"�iJ6�ْ8�ђ�U�:�} ��MݹK^�0�W���Ȁ�Jkɝ��s�<���d������!�꺔����JPC�STZ��Η� ��TO��������?�,�!j[I)�U�*��*!�����ϕ�T��Z��Gk�h\��r�~-�����t��!���M�)�&��v8o��h�,��3:���:yA�AV��KZ|��V�m�mҴ��m�����>�j�$r�$��ؚ\*�aw�<^�R�f� �rOr�O����ˍ-g���14����7=)�*���Ǌ��߾�|�]%��dT'���<%�$�~�|^�y/�У&�ۣ!8O��&YL���J��q��s��g�u�6�r����3�K���� ��0�P�_YՋ���p����O��W��cucc iƱT%S]y���(M��=�!8ZO2(GI���Hgƈ���٨?-�7����/&h)SL�*���2Y޻5M��	�C�h�L����=��'`��-�cZ:�o?h�3��C��E�X=�I���L?g�&'R׋����pm�v���W���Y���}��s8�[Ƨ ���+Lс�[��B�s�Y�ϋ&A�����|^�pJ���}�F< u�ɛ1�hQ9Un��/ ����S�7qDS���jbA�����_Z����9ި4W�����e�T�e�*V.tt�J��n�q�Lg�`��5׮l�\7t�j*%�Tk˄:b9�� ͓)B9���q�ܻk���8L�zF�:�ۉ�~KC�vj���=k�ǻ�����hcF�:h��A���?��T���7+���w���y�;� 
,yⴭ�2Ԋ�oR"L��r�f�ɐ{�`�����|���x���R�O�@��Ez�(�hd� �,HW�ѯ�z��m��r��܂��9�Rs�R醵��r���-��0�%8��}���X.����}�>W��-O
��a�\?��M&Lj�՛B 7�6������*F�c�P,�,Fk�%A�q&��rB- U��҈���ݳ�*
���ǌ��~�����Oq����=3���Y�Iv�@]�r������XU�R���1e��e*F֍��+.	�Ro�ݾ�s/VzPO�B��L��/�Uk�ҒK���ig��1����������a�Q�0.J>U^k[��S�!�^�|����y������}�=R;�����7nɊH�b��S ���u�6 ��8�<%g�����c�3�m�p���I�>�,4�l�w��
�	Iv�I{�A��`���Mx�N/B�����Mɤ�T��I=��@U�TmH�h�0��I�@)MmA��7ͻ3K�iŅ_!�{�1��K��z��)9z���f�kG���15߭'��cu�'�O_����дSmBh۽�P� �@�1���S�$��-�����ryxڤi�;�E�ym�YnBr��2k��^6�g�"��e1} �nrH$�^�y�/��z��#�(R�x�-�k�N��;/-��D*&��9K�]�1��^Մ���F �!���m�H�G�Q=q����;I˧}��dQ(L�sOU�*���{�� �m�Yt ��6U;%�
9:o�M�{�~7�)
�o_L6��G\����~�1��z����	8�����Q�s�UAqNy��Zg�ou�xd���!a�e�?�m[*��@_��y$���!@�9T6T}�,rI��\��̆�5c�����d��Boqg���is�L}���
����o}O�\cy������h`,	+�f]���
�����q�]N�Y�
�<c��c������l+�Ļ	G�o7՜?k��{�u�.wP��{�^J0[��������a}���0�j� <U8{$�\�B z�)��O��s���|�W�������z���u�F����Y�'R��p@/���qPz�1�>���Ӓ�s����o=��g=��]�%��͎�n���G���ĳ��!1]�R����{R��P��i�3Cuh4������t͠�5��	��z��XB���؎!����-�)��.,���{�Y �������6�S�
��%A�|_^I�K$���j:g� ��)���G�缶}�R��Y -�Y�0�7�5N��`ү�}�}]>Y�����Ԧ��@S۽4Y�f�)Ԏc�浘������*�`�O��<�W@񁤵k_}�?���#K�\ �N �5����e8���F�ӎ,҄}3�V�IG�ZK�A��MA�ze:��&���;�ݥ*����C"��h�b)�%�Gl��UR8�{���ޢ͉��ѓ�K�ݾ� (h�a�2���V�$� �o����W�,e�R$i;Rֆ�ݒ��V���Y�q�L�@�� �\i���ah!����<{�0�X�.aJ�"����[�����~�����|��h6>�t�͠��k�8�T+*�E�?`�Y�ʽ�}!|s��n�����>
��<\�l���U��Nг�j�6_Cv�j�����X ���+���*�Հ����	v�;1^��;!D��,?T@]�ռ���>�spw�N́�{����u�Oonv$��_W"���Ixbh�a�m���Фn�*	��N]�4�!������/c-D���i~���郶sr��d;E������U��ߕ&�(@��[�c��O���E��� J���#G�/�c���Lۃ
�<��7�O������[����8;�Z��F9z: ���P~���`���6�5��8:��;�MJ�8����?�k���}7�~�C����;q��WP��k�߹�\�X�[�����+�ױ03�_�^�ʅ��:�_|�=	�:|nZ�\f�Vjn���`�	XL�12��&_ �O�,E_1'�R��K�a� -��z0��؉�j&P��N@ɤH�G�f*�Np���A$��W�r�ݍgy׍�Ý�0󺊂�L�k+��B�M��_k����3^E߫������"�@�ڂ�A��N|��$n�q�Ժ@��	��At֍�]7�v3O�n?� �Iqs���f����Z�fn�8��չx�����C �>��X�[��m�T"Kf�4��T?�/�l��/dI��:���n�_�#6�k��ڛ�'s���t�&u͟u����1k˯1jI\�%��r�-��nBҮҋ�se�*���VȀ9��}�7��q�D�(���v*��3���mu$Lݼ�zQe�L�������`�zO[Z�
Gv�r��� D&p�	��-�'��H1�Ƶ��G(l�˅�������H1����A�^�YYp����s"���@]�c�/SV;(X���[5�vJ#�5��J`�f�ȿ�8���q@���p�����㧀ʽe�c��O�������O�1�Tԭ1�z1P��+J���4sr�7F8�ͦ�X��RPĠv��dH=K�c��A����$��U��z�1��6O������^�ƺ����`����� ]<:��+M��$�ekj�K%�|`��N<�9�HG��]�G���합�? i���~y���n|@�i�gO�L󨸌S�B}��=��>�]ix9������ەB����>J 3�ƳA�pB��m��k���kn~������9��	��I�-�U��n��͞����Q��!�Y��MJ��tt����]��=7��C�-?Z$#)�&)�g��ɒ��0��䒜�!����m0��'�D�F!(i�Nj�"?'��2a���bz�Sy�|^�#Ѽy8U�b��`�$E�E;�7�C�E��0�0���Ȧم��I��O�@���F�Yo���I��?:��@���A��$�����'Y����J�;��t~�8~��E�g�����<��PoM\+ &U�ܜ���Y��&��=��0d�#�Л�4��� p�I[^�۾v�w|��e��^��콘o�w�b&9ڟ�h�4����^�������
	���s,>��i��qR��������GA���3@�����oUn�b5%&�^��J6�j��3�^;�;����NR�9�(���|��f���ُ���K����"�Ğ��	�)�0�B��O����(�ctn��f�9P�������s����֑�ޖ�ٿ	i�(��v~A�b��~��c� |K�@f]I�3�`yK��Ųi�ȗ��o�ύ���*XXf�����av.� (M�b�u�u�[{��ijz��r�"�r�&�*�p���6��4"Z]����Dv��csS�}>����-�ksAݛ�C��x��sZ�e�����c�݈���q��������hhѴ�4�W�->�a7U�5JD�8�R�Km��o��o�v�0D�����d3tIu�L�.����:)���^�X��r�,&�'TU��k.,ؾ���72��SS���p�J�H|�+0Am��!�\k>!=dIĞ��}u,0��{9/�7��Uhl
O�`��ɶ �6Cum���կޏ"GN׾I��\s�3=� `4ڄ(М�X1�M�n&�֖^���#�cP��2"$�{yٿ��tZ��^�1�lŮ�&��i_ r~e�>��i��+8)3w�$R.�~Mt&��� O���8�}�lx�լ��d�iz��0s/N���6��f��u��5��- ،h�=伨ip�$!��#�cZ�iH0�,!k [���n�J��������>�y�M�?�B��s�_����̀��|b�c���ݕ"w��x����w1���i�hݑ���y��s*k�*D��-&����>ݾ4��g��C]륊V��Zxi��
jZP�6�a�[�6._]��j�	JL�J] ��|�ٚ���ժ�.�wڻ��X����NǺ�"���o'�Z^����0Tr��
�I��. J}�"�Y���uIL���ǖ�$(%2��/�!b+�Tf��*�����k�*�4��Л�x�#b�����=��g �M�7�M�3Q��@�Sl��Q���D뫫���/2�8�7�p9�(h��r����xL
��W��"'A+Ƚ�=|�p��m#vu��q�o�S��f`��������~�/���6#'�g%!�c}�o�NW\��(�>.��3��^������5��s�B$:N����4�"��v5�Sf�؁&DP����G�E�zhS�����&~��왪�	?燦��R/�cV��5���B��H�3.����6�����G�[�T��T}t=V��ռ��%O2�Z��[���ǥ�ۜL�H�3���D�(���+�a>o��wB��B�z#J9��脥Y�_�PH�!V=� ��&�;�D�٦}�V�����X���ma���w�1�o����a+ȞB�M�q�	CUo�zɅ��ՠ�[��[f�i�'祓�R��p���룐������|�Hѹ��E���#~��N�Y�j;�@9ڨ�;%t?�����Tck
��D�`[��_���{�+����H6#P'����M�}]II��V���kYߚ��:�df��i 2:7Jd��[f���6oj��5�?���O���Q��z�B<��M����BWx*����ʁF� H�B5�DKa�k7l�qvQ:��߳�^�� ����C��t9K�n�CMH�g��R�|�?@���C�97�%L�F'�V�j�vo-&�uXA�W�T�l\g�����-r����hǘ�-�F(=��ͩ���6/Jm1����ut~���Dx���'N�x^~H��+�������X·D�XP� x�=��tTl�f0j'$�={l�Q�x�K�������^.�56��{*��Tg3� �2������sG>W��["4Q}����.Ǯ��-�aVdt�>�����i��^~����Ս��<�a��Wʞ��{m�����	?�|�Q:W`�T�)Q�ؐ�6X�Bq-�	���\�p�K@9ݿV[^ ��/fy"Gm��}�X)%��:�FE��Sq*V*�>}��Qn���F�)1�#7i�(��"���ԧ7w��=��WR:-���RSqaA7-�\MAT�f����}4�<N`�JJRE�ŏ�N�!)�jx�Y�����a��[��_ע}d�R6��~�"��/�jn1�O��<�).��]� �C�+)P�ڛ%�]�6��Ș�`?��r#�8�HX7���O9u'
��q�Ŋ��
�ER�1CsS������TŅ�y������C;Z��}4�t>4���ݱ���s���FV����qB=Y�4A}��!���������s���ӛy���}�X��ɉ�c���A�ȆT�Oc�@m�f��B��J#li#��Tr҇hk���	�^��23t�$����	%j�����e�0�ъ����c]��1�I(Z�j������di�U~7��h%�F�k�(�������N�����4���N�i1:�>����sned»DJ����+�Ė�Q�_>\����������>2f��x��`��K�������:&���$�f�yuJσn�r���l��\40�����a��T?�G�=�)EF:Ďn��&���c�5�6����� @q�w<u��YY͑R��-g�F�L[l�P��n��p�P	|��\�=�иo(���7EM��"[4��&���֓�a�a�4��ss(H����`��^^����Ղ+U\L�}˧�$u
bM�m8
L��>���N��ѓ���b  M�6vz�7�*������}�BUfU^.������<�41;�'����S4� (�z�3���O�	�c =��A������1lJV�ɕi,��z��	F����<:���Ѣau��ҧs�<���Cx���H�P#=���u�8�v#)�>r;r��ۭ��H��@(��?�=Y#4�}D"c߲gIZ�JT��K�0�%KQ�U���k�6#K%o4��)YG�f2��y����<������|�=���cv�#�����A�]F%�'ڪe���֥�Ȳ���yLt!���V�*,ln�k��Ѷ]K�~�,�:��3 �r�8�J���v�C�a �R�I�ʅ.w,���:�j��*��}��Ĕ�8��	,�LIa������]TW2d����?�%'b�HJ�_�g���x?��I�/�A'F��"P��y��NG{��sC�*�6{����.���t�耀���d��|���v,�8�\*�y�UT�X�s���I˨j�/e<��)�2�ީg�5{&���|���ύZ\��6~�\T��7 ��� )j��޵�������-�>)J�PrLw�����1��녿��I�x�}!��V3ϴ����A����3�)Pt��A�$�>�i�_,x�t��f��9��~c�3z߼�J
��~ C{��T��x����G��t0Q�2�"P�}�x��S���V�9,���; $Pj9,1"%'\��3���g�a�^��X��
�P_獆황�y*�X��|Y��!��s`=N�ÔC��6搵J�9���S�*��� ���z��\i��z�K�f��9'�G*&��~q��:R>��������1�(�Ev!_NU�7O�,6\���w�L(CvY���`(H��!¯�[GE5b�[�f��"3/������y�����>�䭺R�V���˟(f�� �AzA�.���7�~�UR��/�J��`i*�A��I�:��$��>\|��a�#|��V�`��@��Z�$�G�	�c%��(�|t�3D&��ggv봬�����{)�$��l9dg�IT/�>���jx�b�s����B<��]+1�R�M4�PI�V��ɺ5#�L�CH�X�YI�0�xͮ2+RB��{�i�as|	�>+N�g<�ʥ��s1RAH4�D\z�xb��-��eP�=	�	�U��j����P�tF��Ko��E� *�S]n�e%�BH&k-�h�o?�){���|֓��.q[6w�<�I>x���FWd��j�m�D�'�c�$�Ւ�Ŗ0jr�A-��0�)(*V8�W���T������+�,�)V8IH9�_�v�'���F����C&@�����<����hU˖�>�ma��ՒNc@���4�Ȩ��Kg�sx�|�ȼ\�ڂ�J�-��D����Ux!N9bQAbV�s�|��g���N>jl!<��wU����C�My�\�؀����D���ON�h�����r�A{_._n{tF��d�?��T�{������C���;��KH�!$���'������ζI$ģ.�vZL��9^�g�ؗhj�7��y��,��:!����� �`t�É�_]&���O��֪~��_[1<U�{;�������ޢ}�4
��(�5�4I!����S�n��E�,yv�����n��+�R��� x�^Z~18y�$��\(�i>
�
/�e��'N�x�ś}��1^S���bI���F�����|`�O��7r�����>qR!n�����^�S��/<��y�<�/�����
(G]� �y!J�)�/�]Ų����$��͏�����xJ>v�Z��D��t�-F�:�?P���(�:��rߴ@C�L��&@c���� �0���U��
����)�f�u�W-�E[�?�c��z��:�|;"v���t7���׍|���L�/�۳4n�[����ؖ� FK/4���휗뚧.^��D����B@Ҁ�T(>q���w�z-o�G����_�����X���d޲k�ы��v#��F�� ކ�B4}d��,c}X;�}(뵇}�x�RMu��׊�\��|/k���'���oM�0*J�5�HE@��#S�K-s�Wba�A�{����p�xJA]���g�7�����Ӭ�8��*�g�����^,��K�_�8��x���h4�TFR�	ܺ���i�����%�&\�v8@��\g<��w��U�x����͛+y@��D��h�w���0�FVԧ������t,�2ay�y�����U��3{��'Mt������U�8a��Ң��[Qk�&=�)�{����0+� ��[������5��s6"EI"���ҷ��q�%��*n
[�9<B�I��ӂDDR+	���&ҹ��/;R�RD��(������'z�\9�����:������J�h�|`��<�z���͙w�}+-g��X
#�`����j#e��J��C��'*��ld�<k�k%���g��{/3Y��׾j:���HL3+	3;����E�� 1�0����,&�RH`EVU�N����=�S�i0�=�#�+�`cGa�H�������+�yZ����V0�{�k�ۅqM�}l���p��[��L�!��<w���03n)���O �Vm�5����������ϓ˪�Jn�>E�Iim�i?�9���4�Ec���
���J"ot"ɀ��7(�zۻV��2����	ѶӨ�@rя�6=��$zWp+���.����!��6X��S���gn�ѱP����~aD'�`o>BpXQ=�Xo�DAѡS�*TV�(ab�I4MpSG��*({��X�˽Xv�I�TH�/�(E8W�䑀�x'�1�5y���w�ҽ�B�а�~�J�BO���ڋV�͙��e{wF�,ǳZ`m�(��SoGm}�
z< _t�C�嗾u���4��텱���������:����L�_��)��>�r����& D�~�l縉�,���U^�����	6*U��I�=��W�9�=q��8���ɟ0B�l��	��b�ď�T��zW��s��EF��qG~]>��k�4��oSq�2�gl�+n����Ƿ}Q�<�Y}Qy>q��t7C�n07$��ܰ��˳�3�L����7*4H؏Uy��mf�o|���U��P([��:<�h�N��⛃�Wa��!������rB�B!��������31�a�"� �;�½r�8�tM���/��&�Vy�O�Q������^ |���տ�)�~�u��C������"S���n�{����e�D�z'��Y����r��N; -����h��8LH���Iƾ~��A 6��~)_�c�Դ,;��b'm�M���ph>�ƫ���L�M�eR��J�F��=�,dV��*���Q�^䘳���Q��krɕ��=������o7���}�|�txA����끯u
��=�����?5��jq���3�������+���i���HU!�O�H��K������J*�m��CHb)0�bj�X�	Y��iL��.���z��Owny|�w}����j���K>����(q�,U�s�:�[�Ev��m#G	�ߎj/q���p�y|���&N�p��3�}4�v80�	1��;��Y�آȷ�ϡ޷K#&!�Q Yt`}$�ki���.�6XhE��`� TAlƄ�����3����<�P������������+s���1_.\b%��!�d�j��?!I��`�P�Ć�G�XMN�$�
6�1��#ʮ|�x	�կ4�/�'��иf%�ؚ|�Wt��S�\�Yr�#�\!tB�,�a����h����>c��҄�n�#Jz��
B��]*oxN��v��R�*�dӌ9CK!�
�s�Zzt�F{�;�G{��3B?�#�g�\�8��+*М�鍆
���r�bL�f�����H���-dt�v� ���p�K8x'
����ƞr[�xQ��EQS�o�i����B�¸=�-����6����sͤ �{>�=蝒{�j�j�� �����El7#��0�ⱏ�U���|Sy�����Z�-v���P�T��2V?��9�Q�����i�x�+�|0:�@�=��}�u�[��ȁd�/��e,)��Del�H6����n�&eY
Tg)�P%+�<bP��T���1Yv�X4ah��q�=���H��+Y�Ǎ�)cnu*гfm!l���q&�5��c<"!��.?HI	�я���]!��@�l�Sȇ����݆Oe�������ѹ�h�����~=8�듯BnW�
�?,2{��j(��+�����ߧD%�>X�'"QNA
��U<�?�}��0">ڻ=AnZ�1��..�<�,b��e�TbS�d�%�sp����@���w��e7�B���l��U_��V5���V�\��#\�c�d@.	;�(>2_Y.Ҽ�ԭu^����ܿZ��yoYҵb�0���b�3��UR�h�U���u�˰�L�c1W�#��@�f2f�[�;G%�����tE���j$4��r_�L���1�n�u����7�Vq�z�h`a� ��O/_O��B��ߠ)�I���1��?�2g	�m�?����T=+k���FФ�w0:FAQ@R)�x�)�^-�/Z��p)sv���X��9��Gop���Y�n>;��R����`�H
@|�� t�}��D	7�\�����; ���?4�JC�Q�F�;%x�;$����̚('M������>G�m�r���n?�7����G�<��$S�QYm��z�S��Fs����>�)8�k!��n��r�u�wnJ�F���� k����1}����^�'&%=
��C��d��n��%���~�x8G��w���v�X�A��/}~�޹'�b����s�o���H�� O�����߯�K���j���$���^A�<�#��lbz�c�k��'"s��!;4�H/�a�Zy�n}���G�/�R�:�t3YL���y��{��F�����5�r�>r�Ҭ�|;o�o���<�����l+^	%L.�4B��ôʝw8C�ZՉ�[l��%3^B�H k�B�r%Ê�����u�y��Z�{�� ,�|���j�昉G���W/��ɑ����A �m|d���]�b�0��
/jb���i4ѱ�U�B�]���L31����\�J��T�u/�,�YI�k9[����k����Åh�=�z3T�q�"|J��Ay�rv��Յ�&wЫ��Vo}�p%^����\��� i��"zZF*�,s����-S�t�����k���Yq�%������0W���J�E����й���`����zӘ��U:S��A(!�?N1� 6��%A�N�&YuǍ�t�+�B���)`�2�
�_��i�s<��'S����FH0��&��������^�}�ף�+���?P��\�#K����Z�
�P֡1�KS#��K[���C������cM�K��¼�>5�I�=
�\�� >�g��[�c�K���qa��W����=�~��m���u�����̈���܏���j�Cq��N���nh�n���״���ZnU:���V�)8�I��ݍ��1�թ��k�	�=2#c��������S-{���Q����JW������Hna��qʮ��Z��\!���QNJ� 7~����;�*��y���YwѲG��������;&�^
2�gT��#]���n?����`�Е����&5� 7);�ќ�݄��=ƃ$�j*�q�U��p\��w�[X�6�i&�v Hܰ�T����K�u^ĵ�!G��O�E�f����괬<�*�y�xʑ�"yߩ�c11��Nf�_9�9�kr��UD$�]s���$�~�Qh�r
t̛,-�8�I�R��eu�4��!��"���  �_���bV≠�ԅGk�Y�8����$��!��o���W�;��v�[���M�tޔ8��)��܅�o�S�\�g�x95��45�s�:v0{�������Э�n��ҥ0�����gqh�����֥��>5�C�)j�4C'
:��H*Zԫ!��=�\��0m�K�k�-� ����݁\�w5�*�Eg�E��п�k�{�Uv}�ْ."S!E������:^�&���S��'�q�v��&�]arR� �0fs��f�����ڍ拘1_���Ctz����r�����Ų��p�1�bZ� &�DY~��^��f��4���I
���V��Z�uL�a+�^݊6�k�)jT#��ã�v�T	�q��m�
9����F|T$����	%�H!�+�����Y�Ftm^ ���d*Ე���g�V�ͽ８t.��m �o�ˡ��?�䎣ce��eU��;� .k�b}ׄ�~_Q#�rCxBf蝅�,j5�	�sP��SH��N��l��Ue�R&]��$��꿡Opn���N+A�[6�P�� P��<�r\��*��B�����K(��'�B��d�/7#$��Yv�Τ�J��Uhؙ���k�.AE'�4��_Π�=i��3d!c̊��V�0��S���lGM3��A�D}��	�f����+������`�=�]&7 � =��d���&'$��$V6.�pҹp(��$]Y�P>���f�%��7��)�$
U���,������fW��YR���U��^M�	05c��+���~��rK�?�f �,��KeK��̛�m��Η�J &�$m�쎳�����s?�?��B1�*�?~9X�ɢ��i�����0�K��	��X;���}݇g>N�V���<�ex�%�r��3?�}�����w�ɹ�N�^���w�H33Ա���f��j�cW�l8k~x�<�(���H4�8���.�4��>���r����O����0+T�`��q޿���`k���7�)4�V/�<ֱ=k_=�q���/��(�X�,��խ׶�����pv�=�m�zVN���n;�R���^K�k�x�7�"�>L 換�
��������i��b�Rѭ��&8ek`r�ɦ�`��MH���6�*HG� �&��x���	k�8.�<�N�13�Cg����r��^�NH�ЎV^F���3	�1G�o�y�b���#g��H?-�r&��Ġ�� �/?'4A߫��/�uO�sr���Vy5�!�� �$�l�5��<�W>�Pgz"�H� ���1^�ڛ~0� g@�?�hd�p��50��,Y�Ԧ�9��<C��|�Ժ��{��h��`-����}՟�I'��{L���/��?R�G����$�$����o����	y�7�tg���=�	�)`}�E�4K�%�ի�7ߘ�LC-Q��,XRuj�?��b�P����~�|9m�S�SRpaTQ�W��Gٲ���=�+\�*r�C*t)�`�RbK���T��}g�.R�����gI���e�}r���Ĕ|O$^�-���0�7���(G�'ū�}�c�'~\~<�Atn��)�f��yS%��ɋo�s���k�v�6�h��ê䓄єH�K�_r�F,�	���͵mhV1^�:�4~=�L[���,/�p^�b`�F�A�mk�Ǭun� ����ƔŵM��*�g���룛/^����a
B_�M6z ���>0�#-gyC���0��;➄ ^r��+���1�A�B�T$"ބq��޷��ӼC��%yIz;����,f~���%NF�J���M��M�ƙ�)H��O���L�m�c�_ZM�~H�����r�������V�-�����M�&+������AB��ўO!|0�ssB6�b�$3�~�Y�V�1�ϑ�O�6�ܫ�	Y�}�!����_b�5��%�N��^�R)���D�qaV�"H��;m�(�P�[��q��G��8Z&��Ղ[R��v��`%#P�
�r��\�.�`���C�Q�`�QK�2��kv�9�Awv�;������TTV���0{_0h9��τ�� |C4�҉��r�l�@8�k�̗vh*�-�^�����\�]=������S�{.y0x���d��3Q��yNr����2w�]�2v�;:Q���+�E�;���(��#�B�Te���߂f�f�U.V�����13�A�wKû�@��ڀ��75[&��_?*<z鹞�
�6�܍����'g�N;�Pm�4������
6�N��bA1���Y&���=�����~�h�ɩ�<�Le��,�!�,2C�NB0I|�46��.��4��d}���-��ܠ���o*�`�n�P�n��Q�i�H�`z��1!���[1��W��T�4�]�=��;�^.`�$�� '���Ꮇc!�g]���s�٬���z^�y����gx[b&Qw9�hw� v�1_P�z/j�}E�(�K� /�"1�v0_�9ʵD�k��^��6
LqaO� �n��f7q��)�(R��E*��caDY����X�8��~1��6����tU��a�P�r�ΎW'��I����q#�vJ���W~�A�OW�q�����0����E)f�׀H�O��e�݄�g��k8�����h&�(�]�5?����Aj����R��e7��H�˭e.��,�ejN<��ጺf�v�>�,�1�Cbf��4Q����2=ڣ>��8����c��Af������[�(��v�\��Lf��8���o��~���Z�s`1�$&��~�C�
�S��<*P��Ǜ�"�I�C�P�vF]��ѥ7�<J����啼�I�q-�(5��D�V�����o���?N��nR��/,SS��̖V��S[k&�l�S�L�����
i�z=�;�I�s�${~���RH��sŃlo�7�̓��UG���1+�B9R�����v�B���>���{�Y�qz3/
� ��o`���u���!�6Uk�g��cK��2���Џ����t^�̾���8�(ł� |�A��к����Â��И�"7�� �y��,\R!��,g+���q&���U�i6�� ��ؚ�B��U�OUg��-S9/�I��? Ӕ��[Z�U`o�W~H�L>��H�?e�T<Kjꔳ-�<��K��1���D�n7|�iÃ����c�����C(h����6*�~�fyB>c�qr��r"�sP�0��cg����^\���{�5U��)�E,��?�N��!kL���E��Br�lG ��t�>Ž}!�=���ɚ�!2��p���R�^�Ƀ"y��M�^ԙ٥�CȾ6=VLi~�?����T��q�v���[�/�V��y"T4.T�{j�Il�;
��~�621��1	�<���U�`l� �4ɇw݆��!����u.�Y�Q��A d/���>�ל�㨞ó��#c�xxKD��-�2Q��
�lk�})>�,(���U}�2�Y�:�ԛ[ze��CH96V���.�AΛu�;�&`R]f�ǌ7�Y�n��y�Dx�H�n+s�V7W*�g�j��C��)��Yu�����f
�yL0��e��?ɞ�x[�������	�uŴ�O}_Xz
U�xn��j�����*c���+d˚�����N���,����,�a�v<�c��r=)?F��D��\&]Ô�S$`?Z%;4��C�u��0ˋ��^����O�j��u�y��[�0�]�F3���n��*����YF��w�[]gpRX`!�Mm��E�_�^m��1$G�݁�+�!�J:5�tfە�����H?�|et�B�m[[~�[�|\����q>�1�eTA�.@COh�7��H&y$B��wT�dْ vC@lbM�sCLY�c�򾸃�z A�L�n�(�R�n��tg�]hc^C��S m��B_�V�:�F��ʩ�P��#w������`�L���u����n6�ܫP�/~dx��DVm� �-�S6��u��	^G���x)M�����#��ONU��B`�#z5�o�m4�:(���#gi��n<���t�+�9-��s>v��_���X8�t������~������������`�E*��If�oZ@ֹ��G�_IS�d���?��)팭]�`4�i�FlLC����m<��+�0%�]+�t8��]HP��)������v�v�k��I�[�f��9́���Y���]5s֑R3u�S��P�M `�������l��BG��K�9�la�RQ\��gaObi��]~��t 3؍�e$դ�3]�$����rS
I�|ɲ]+lD G��yF�������(�!W1E�Bsa�i��|lXw2�k�9��m�=F't���)��p<�!����t�-���|s�/u�n�� [�]6/�-��8�!�������`Kx" ��p�S��8�/(]�M�Oy����a|u�\�=a��Ͼת(��WC�q3N{�Ե���鼔��?�~���Q��w�w��v���G�u�-7my�|�Zދ{���J�A.`$�0����^S�彃��!�ͼE�r29P�S�g�ԧ�3Ղ�����)���,�9\h��'չ<P�����Xv��_+�4�_������X��z��ɋ��)��J|�/^�w�nhυ^���;,����}��N�p�]u�znt��w���CH�&�HZU&�n��t~DU*����II�9j>���Zy3�U |� ��e29m�p���� ���\�p���ꡏy��\�0��м�a(�3T.�q�8�a_��� �?'�2@������&���ms#�a��u��Ƹ���P�b��l������ǅ��V\,26�(ꥊ�z �A��9��X�5�F�g�^�E%e|��\�*r=�JJz��G�Qi>��n��H�!D�g�M؍�[���⥈��|��bLK_��25Q[��pU
6�W�����C}�B��Ω�64M
��S꿎��ڌ�H%`�RIKǼm�bo��˾���9� 1�O��Ue��k��R;L�CHI�!D׬�t���g��2�o�&��[P�C�"q3�.7ܽ����]� y�p"��<  �<Zr�hE�]���YT�㏤����Rn��҇����g��ml�*�l�%�"������b4xd�Z�'�NM�]��a�%�j� �bL����|�g�y��?�q��O}�t����ph Ղ������7�ÏCW���%V��nF ��t�ko6'^���4��^��hC(�uO�D��\�;�ۣ�V6��J�5���ǈ���cD�<!k���Ȟ��X�Z��1��mɘ�B8��#=����,�*]�r�����C�%������9�<�4l�~����L��b�5ɚR�L6�i�~7H!���F�e�G\�q��ھh�Y:���D�D����I�b�}�hsN'C��Yҁ��/���QДGJ*y��������6��:]��Vm�{�?�z���F���fZ�`�G?F�rv�-s��Q6�1+��+<>A@:*B�o�6*�g��Q�b3.Ծ�/'�6� �I���訲Ύ5V0�}k#0T�L�C��Y�-���V�5�#��ۤz�u��:@��ﮣ��_�^Y[;NeuqY~]����dXa�L�W��W{�i`5�`����n/�M=+���������{��Do�I�&R�N�HIL.iD��0��D_��Y�tvI2���V2:0�7����ϖ	x��$E��]�bB�2�#���z�,��������V#���I��)/�bW�m���)?YJ�":H��d�����O��]Y5Ӟ�6�����W6��������W�y�O�D[p���%�E�Df���`>@��i����vk�E7JH��������q��se��u�.�(�K*�;;=lL 5u̬Da�S7�{�c�T��LpB��T���w�K耱��a��kQ5-����`��{�6� '�0c��=V6�x��f����	]K6s�1�Q/�G�#!��m��z�5�V���_�drR
�����O��O�-��2��%�o�6B4�(�ѧp�eyn�f��~��w�唬y�
��_.�y�i��&���k.��n�i$"�3;]_+��Ԭ_n_��l5Ҕ����l�dl��� ����1P���$��(G���!�ۮ0+�Q7?��A
�}��~�6�buF3)��c���/%U�q�o4��+,	���R����#e�M���O��P���|���6ػ _/�7@���߷��}5�����6��J�������u�W	uu�h-�bM7t��fV�(����L���`���J׃A�8��dV�D<ɮ�v7�"�n�*�V3�.��_;����_0�뤸IOb�����!�7���v|VR���G�%e��.~ȈZ*L(͑v�C�hng�L������-�!p�XA�|���OIe+瓿�yQ�y�����*�t>Z�}/?���p�O��n�"8�6��XT>i���?���D|3T,�~K�݃�]k�<m�����+t"��#?���{�9ť�c�ZL�qo�苘0����$h];zBڭf141V���Hڷ'D3"����G$��pktEɱz��+���TyG>��9j,���~^���*i{O��$x����J�Q�y�*�[X%bc� ���Ş�=K���X��姚�Xs�x�/��a{=�`.%�ػ�*(%jĖF�L5'��둪,�]��M��tm���<}��%�e�������_]��qp.p�^DB�/��e��� ��`�@�2 8-���3�<���ג�_�|[�b�h �`��k��{�:��-B5I�����ph����>�cv�u�G}u�LI�2�����	WL�i]�Q^_򑯄�������3�t����%�,����F�R)�k&I �_�YXC�vk�$��(�+ ��8��@��d�Fq�+��|���*��A��׵���T5X�x�ʿ�z�,%t�W!�[�v ��΅41�5m���ƹ�#+�r�	��uۯ��:(pT��#�^tbg�)Y��� �~hr,5�R����Q�l'!�`�%I�2CM֒G���BRx1���L9+x7�V\?rN*�lzR���g���P�J#UZ��>�?E<��iS�lTW:�&�Xu3>����(���� |�+���JI���V��(k5|��mN6�>DL��qR�Ǝ�����(�F�i͜�r�a��N�]�
��R�!;�^t:���*�%z�����(��+b������ ���b�����g���{��d���1��$�h�&�Qԕr���]�}dS:cl�tb��+۰�B����M�"T�r|�<�R#ܳ2 �^��Y��Nq�L� |�#�F�@!Q� �!�4 ��};�{En��r����k����X]�~��*`����ۋ߽�.yJ��x�Y4Ϋ-��U��=��*&dWs?��0���fF1`j0��i)�ޗ��n��Zh�U
rp�������佤�b^�u&�������n[���yN�stM�K�M��A`S?��<UlX�4yx�B����t.�:k��e�������WBt�-l��5m����|�r>���M��L������U����7�����l�:�C�3f��[�	���@P�v��׬j%����Ec���Ɛx�1p��������ЛNg�g�K'���2����f��:��J�e+b��s�g>�:C��"��}�MW,�+��b�M�7\t�X�������/#��]Oo�VA�BF��X8-�j#w��?�F1��M�Yai��,V4r]M\�ei�婼"	T�ό����TtN�_�������۾헆.	� ������4a�`��m���yb�W��G�@<<&��k�og��s�V��,Ǔb  )ȕ��5-�2Gk�K����Yw�l��S�f0�������T�q�<���<����Q�s��̝*�+{J�ģN=ab��僟\�e��6<��2{`ф�r�2K���eVQLyմO���mt5��}��B�<�k�g���!Q����A|�EYۼ����S�w&1����2B���5﫪Ǆ��%Q�΢岑�n.����|}r,<�����1����)3H1�uj	�e^��k5��rb���#P2`�y�D�j܏Í�S�����A�"h�`�����K��Sy�~8���{�,�!d�g���{q7�T;�+�Oblu��U��~�R�����t�$�`ڿu�A@ċ�*�r��q��RW�7�ȳ����%���Ew%����� Vu3�`�J�v�J�
�-*��3�}������ϫwe���P�N���8����jܙm����=�H'�"���]��߱����[.N���?
��D&������Ȼ^%r2z�.��7$�#�`YlyD��|���z��8� �EqLCp�ϴ�}�BY��j�Nn6�J�`�(���>�Y&JlP*�)��
���)I�tp�P�d����ܞ�G���Q[S��!D�N.)�ɜ)�tӯ����p�D*�=I�)���Bh�W�k�Fl?4�:l?��[��:zDI�����N܆��G����Y��_�+��x�|;S$���$�kD��#@���>?��"�;��?�q���}sݎ�7���N�8�k���j���D�ؒv���S@B�1����6a}QbV�Y�h�\ b�G_�Ppޡ��Ey^��Ԝ����F����������^Y(��mr��*=��H�c��Udu�>ي|��i`C'�c
2!��c�FIw��n����\���&�!R��N ���9�{�J����(�}D7��<)򶬞��v�����0��6�{�[�t(؆α���Ց�Ըw��c˹���,����`ݬd*�/e�>��d)��Hx��W��7ł�}�M|�׉O�jhAC庽,��rH�Ȭ�}br�bC!N�1��܃��TB�!��� ��&�a7�l�N�TU7Iv�����{<|�ӂϣ��7ƚ
��B�� l��G���m�zC�j=a!��E,Lx�x�1m�Ӈ��担ׇ��'��2�?��o����y�'�FbDr�hwV�;ަbp��Q2�#�s�̌����u)� �?�c奯��7֞�ް�mf�n�z�G-���w���8X�uW������+�F���[3
�	��`�����,#�6�9�r�g!
$ܷm�_d��L��)�� �'��s+>���lƙD���߾���OY�e�.E�F2�"?��K�IV��?��>�z|E�C���v#�Y	���[g��]��t���3����j)�g��	(S�8�W����̎�D$�CH50�^���Z?��ޖ�+��:���0]���r,���N����Ou86U��%{(��i�E��wᰏ��%��
����.o��^��*�Uj�ηE���Gw�=T�&:9kY�=�e;�+n��*�r5���Q�+��r,l�#��K%3������t�$������-8����bS�nl���B�^+���@*� ���ݯ��i������'�b̀�,ڏ�L�\Զ���"L�me=c�&�VP����;�G�ڄ���h|"�1�+�]
�y�.�wz^ٳ��LrB]�JJ:Bqs.����~uފ�r"&EJ1"��뺋����]U����-��1"Y��H4����ӎX����=�]8�q���>+�T�A�Yګ�W��eãjh�1l/���@>�n@k��%"�b�����W�v��.CeE���4.�o�����)S�e�^8�y��?�9�@�ͮ���ߍ˾�cc9E�C�����N��=�*:~:�Et��8&�����C���vq;�v��5���t�V��>4�����|��.�@F��e��=��{�O���|~�CK��jrQ��s�8��q�R$�r�34f����q��&� �5��5��KP%� Td%}���(�O ��;?�?��\���&B����
��eNw�־�� h0둛���Q�_��"�Z;�;�=b[jL�2�V�ow�X��y��	�^<a�lK��G��/'��ֈ��^U��9no:���s�Cռ�Z	�	��,qX�D?69H��{�`Z��i���0����1���`0��}��'��B�OT��u���U�gZ��J�ۿ��k|W�)�[J&��A����)�������-h4{~p���W?q��HB�9����vT($���g���Ht�7n"���b�3���D����Rk����芓{ �t�nб��Kɨґf1��x�	�HA�K4��x�h���� ysp�nK5�L<���4}���+�Γ��F ���I�1��y��N��bz؂Hc_+ު��)7�'5���䰕��P��rO�V+�5�!���mx���L��u����]Ӓ�����RY�Z{�~����Nn�wg2_Z��T&�$IX��N8��Z�]����OKF�Q$�q:��/?�/C�_2��!�P��� OD�m������͜�L!�ek�' �	�9jXjg��a�"�BZ�@����	 ��9;s��U$��UB�_d�Jb�.�Ƃ����(%-E���7��;�D������_<���I�'>�U�QU���Rc�(�#M�%�]����v�������2S�ۉ-�&�c��g�`�*� s��E�'ۢ����(�KE�����\U�ٲy�M�uk���5m���b�S�7u�褸��J1�=�͋�ՠ.f��Os�s��o��)9�t��*5[��GL僄���r�`&(j
|�yq�ycG���{��� %^6�+��B�"4��0�L ����>����ȴe��c���X3�w�Rmk���`�I��ҙf�`齻�O��9W�5� 6e�����%=o�~�[0L1~�QQ��7�/}�R�����{�b:A��De��Df@�Bβ)�}�F�d��I����7����a�lQ�~ʏ�cv�N�I`�+P��^#�e7���J�9�7n��L
Ƨ�V�ee~�R��]'�~�`"�@����f��_�%��^�b�ȭ�y��˾ 
�{D�~���O�՝�{y�4���L@�����X�gѝ1&2��T[B$ "Ȣ�	��0�?�Tb�-	xn��~~&.x���?�C\���x��d�S`^�X�6��B�	[�n�{�xv�S���W�hBV���}�Y�2����b��q�"�U����<������ LԱk�5�0�KƢ[kY[��.�S�]|�c]*�-_9�5*�m�j ?�P8� ����2�[����A����l1��G��R���p1�ݳ�����+�K*��Ws˽ƭ�pKM���ǋ�ij�d�5�k;��'�d����k�Y����V�%n#��R����C�E.`%�w/������s���7Ѽ%̽��e
�;�jH]\n��\cm�pu��-¸خwF�Q4	��3b�e���A��UՋ��4� '�⌑��m��եڲ�r�>� �����!B�hE��s7�P�<{�)�8�a"�	�؅�]�>WtS�fQ�%��	Y��)�CϒZ�/���NSPBCE��Ś��ھ*���ل<@w��0d� �7�(a�O�&�^���	���o/�D^k���3R[J�_n>�ĸz�d�S�J;���E�yHf��.�zj�|��և|�Z�vjE��H��P���%ڳͼ؂�!Oƽ����Ȼ
�"ٰEwL���U����n����QLM��i[�{�cj���L$��m���U�8R�,�-~/~������A�!�[%G��#��+�r�i7�b9J0p���|DR��~�'GF����P?��6����⺊��9�q�tt���U�3�#r�'D �z=�l�9N>E�	`���D��� ��R�b���`���x�q`q�	y�G����`L��	�w�,l���L��
�O�
��3�V�}% ��s�vr��ۘ*�	��N>��;���o��.� ��/Jo2T�,��r�����K�=T2r�Y��D�>�F lL��鋪���	�؝���
���7{�x֝�_����;��)W��`J6�;ߪ��U.ϹQi[2��㳒����V��	��&/����H9f�c�D�r�IENq��u6��:Ϯ,vʱ\��^3����(^90bj��`唗r`���-�����q�7��͒��Lw## �嶩ug/8��P���L8t�"�f�<!T)*K �'�aQ�=wLƣp�\4�*_�:7Ƶg���Nn1,D��fĵ���şBl+\f�=�7�MWdDW����x>X���<^��j`��wg������W�4��&3��J �o$qk##r»��@�4��Mt��A��m��MmW���)Sҏ�Q�V]�xҏr��N!�u���>�P�&kc6��:�2��fjz����b'oޫ�!�"AE�B��ai�{ �^��|��hL����hU}�&;���f�K5��
~�j:(ΧA��ioj�?�����2������`c)��iE�~���>SvRݷ[��\!ADe8	s�Ýp�]��^��74�� ��)z�Ƒy�1:��)_d5	�tE�%)|l/�Rb����O�Rl��Dz���X$��P����e09�G���^
�I���thei��]<�&�.��a�>�z��F���W|y�v���*	P�W�҂�u�"l)}i�\l[/$d��Ԗ��hN�X�ϟ1V�ݞ����u]^#k�k�� ���6LH}tۓx�����2�=����>�-|���^�l�K�%�v�ܸ�ɾ��J2��ڵ��Ng��H&Tpi�t��5|#8d�S{� �$gQ?4
��	xة͡Ҥy?0�*��(��P�x�~�#�3k.�W�ʕb�΂ ��	�`���cr���2Vy�����?��I�����v�!0�z�n�4j3��p�b���.�{�ia�z=�S�U���Mꕜ�E�̗WY�M{��#�-�p��M�.KӋ���uw������*F���:�����D��r���tV!ȑ�m5�˽�9��za�U8̳�R�.��J�]6a������q;�đ�4�Uh�T6{!=m_�������<R ���o(ʪ�ּ^#�e�] -����[�g�N���G�[/E;P��{@6'�/����ؤC�_yj=��Ns���z�m�+<��<.b[��%?T+n, ��ݧ٪\C�n��N?�X6#LK�&U¥���7O�gL���"�e�$v��o��%S���Fj�}{��U��WW��o�q�ܛ�ɺMzi(δ��'��JaX����X�\�*c��!,#���!,����[�t�Ƃ��a~�Y)^������{��>8�hx��x�l	�˸��ͭ�D �����Zl���-��;+�=c:\J� H 8K�Q���2/֙�]�T��ܠJ�L^�Nr�/��0F����;�	� r�Mq�Wo���B�.|�Y�k�@�(p�&���/�F!��XR�f"S��BHf�!�F4�)����`0@O��'�V�WP���ĥ��$��s|�p"���%@P��Uj��c��VN��ܤT�w�X�q=����a�STY�B�G}^�h�� ٓ������P��[�,Vw��u���z�H�����m2�`�� �1���h�P�~��RŬ����(v!�y!��6&�B���m�-T���M�&���> z���gB�I��f�% H���^հo���i'佬�$��> �x�zJ�S�X��۴�����R{o���V,��(&�+�E=p ��6#�K\ɿ��5G��+R�]�����t���r�)*k�A����_j�U�`���3�δ�1�����y��Pލ���g+�#څ�����r^���
�n�[a�>%3ʁ���<̩?��h5��@j}Nz(Z�6"���^�`����<�S|���҄����ft6V7����I|��xNna�@(.t��z͝�)n�Y��*F�xI=����]�},�=�#\���on�LD�����	��,�:�W;�>{��Ȝ؅<;+����N��D=�k��x7�OXy�=2~J�MD�o�Jt������8:�jkUzh��݌j@�H�Y�͵�)7>"��O&�h��6��,��Q���n�D�M#��!B_X<.TƜtv�sy�a<��w~����N|����c�x�'��� �d�#���ї���R�����dH��[��b���6]alF�0�{M�P��]0z<��:���5����̊CoI�Ў=�h�����=I�z�E4kGX�a�9������n��5���?3�Q����YB�y�#�(&*�\+��'��/RAxz���$���L�PK   �R�T��K� 	� /   images/cd1eebff-8d4c-4172-8358-6f93b12ef793.png V@���PNG

   IHDR  }  �   ���    IDATx��ߏ$�u&��s̬���_"��hDZn��� �o۲��4���/k���a�w~�_�I�a�G?�����&�ZY��"���RI\��a�L�Ȫʌ������U]]���=�3��}+3�Fܸy���q	l��l�����k�?,N;�|��8�l����R�:}쾺w���=Q��O�A+�{�p��ݍ������W�컗o���4�A���Ʊ66VE	3�3�1 ��L���|bwG�� ����E�Mk��`�c�T�fK�<k;���. ��p�<!�ݱ~3M��5�����6 $�� �Il-1��h4�a7��.��$��)�ԕ $����9A�:0� ���Ա�x�֭��#ߍ6X���`�VA�e\�v:���W��l����O��TCn��>�2r�������yf�/�i绺�G7n�:pف7�x��4�8����W��*� p㪝<���ת[��������1p]q�j��]����󋴽���X^G�S�G]�X�}wkw�
9�nW��n�k�/ �_�s��?����l��2� |0����h~{��v�Wf_��ӿtܸj��օ�D��Cuk���a�l�����f\���X�{�u��?�[;��/L;���_����z5`�Ez�ƴh���K�H'wk�����bq� �`w¹=��k���=%M-����|��&�k׭#b�iD `㎪v� x4�̈��e]s"	�睙���6hѨb֜Ț�4' m���d�*�Â�ĬaȊ(pqA�HJ*Mt�5���B�f��^�֑��X�Ξ�� �)�8�bĉ��OeѶ����,���[7o���y6���!}l��5��=�ғ�a�m�}���)��bw������-(�)]�-�i�`5O��#	�[�)�w R{��;"4<� �6Y�������wp/D ��˽�ד�t��v�Ȓ�R� f��(��Y\�JnJ�.@�EʒR�q��C �� �$Χ��� ���vN��Q2�7L�0ClG6�����	�g��{��>_Mp�s���1kZ����m�J��I���%�� P�HM�XP��5�&��BV�e���u�6k8f�ց_�T�u6��*�͕@]��
��4Kpk2@L�LFU��Ɠ����Z�"8 t�� ��YNۉ���'GSG�G�=O4����f��� ���i&sj<�mQ�q�g"��a�� i!\+tЃ��`�Ľ�`����j�W�ա�\ p6�yE(*1��2���0	@Y�j�q��gU<;H��nr �܌HX��p
�.��s���$vD�E���;XjZ���L��Kp�2A��T�X$����@�DN�Ⱦ �]u�ZR��f֌����o/��ݽ���p����|�!}l�cUm:������y�"���M�tA�BKVg �v��dm�Q�	 (Ufi�j$k��y���q�j�$!x�����.$�<�@��N��I�R�Y���C�:��Db����8J�kEu��"ޒ�*�N
��)~��-u0��F�+}. ��%q#� A
 -w�<">`UE�zb�j0��J �K�	�]�,��m� 0� ���8����$1֛�L#�*y)��Lr
�6��+ `/����� �������o3g*���K��4j���fdB,p1#6@�0Aۗ�3y&
�uq3�A������ȉ��!3w�35�fX�laf�1�HJ�89( D�D,�Np0*7�	�
^8�1S�1�_��Զ`6��#0܍�����O;�����[�Z(�`"8;� b��#r L��;�`�`q5��s7V�����sbe��`'r�	�N쀁�H]�D��0�3�3��RZ�؅@D�09��	�n��@p����F7��0� ܏���Cs��2��R7���_Q������_�o�����gkU�6xHlH��k�P������u\[�e�n ��#��l6��t��z��~�����eH���l|)H��/��t���\�[��Vs�q��W��v߸���׿Y���y��W�~�P����E1{e6��f^U��������鬻��� ���Oo������ʕo����On�� ���6�{�h�s�;�=':�;0 i�"�Q�u��ig�Uv�ˣ<ˉC�jO��խ�LRp���dZ��!�LZn�"�V)զd1RmYTr�,�� b䦤��X3s��������,,Ɉ �F�E�č��؜� 5�T�M��Ɉ؉p7B�.�Q`!� pa 7�Hԩ� R����ȸa�ƍ����Bd��I 8ca�#n��HU�*�km��NRiCw(��``("mXi˴���fi�Nn��d�7�12KHn�q<y[�@��n�R�9�<.�.�Z���ͣ�	1س�XXA�P��!����ȁTc�P@ b1��"Av�����Y�FB!!�`���6S7 �X21��3`�&8���� �r�@@V%*���ЇBDH�F �b�;�PJ��>��/ڗ��9/��{� ��X���D������%]~��%���BVEd9��&�����Y�DC@D`n���B������!�CX��>�Q����]��n�q@���~��27�aC��U\�����/�'��ݳ�싴XܦU_���6��>���C�����Rj�mƥb� �[e��>���{����lF7o~K�\�'r�������7?� ��Po �}���-��Ɏ5{����3�9�:z߫��l?���7��x�Σm ���6 pIw����kw�_�A�\�Ej_ݧ����+W~"7_�m�߄��7��ۣ���������ݶ�"\
5�٪�ȉ�N�|���G�Ż���&�CUo�t2��UK<χbR�w�I�B��#
 �/Q��(��S�J;��[ud ����/0Y�^Ea ��H͹jY�MI` �$�Y���)1��D�b�\A��8���ڲ����K��Y���q���q��Dn��T	lDfS׼��;3�AA� 2搌� �n@�n�pb���s�ى�����48,�A�M܉��9iMd�
n��V�1p�C�e^'"q��9P��R?/ܼb��j$��H8�~:P���{����rm� ة�O�;ء�B�@M���RO&�0d�I�	 ���ݝ�(lD���{S�9 �Q육؁�2�A��L`�
��s ��[���v���,�O�L0U���
���0@������(�
f'߫����0QO��i#��`�c� 1AXp8?@�����f�5"Z!�=��^i#�e�$h��| g�*��,�\U%x6dS1BX`pXV�	n��@� f�!<��렙A!�0xT��9�Ӻ��o�U���|�'����_�c�΁�&黶�\�t/��~�3����+s���6�?���72��?`�8ׯ��.��w��]��b ��4dO�J�/K�����ɓ�ҜbyJs��?��v�"K����2����fʾȦ�8�X��b䣼4���#�"�(Q�"S�r���X�`ɫ�7�,�w�u�h��� 8|���H���F�)%WH�!���� RU�P	{  TIn�¹�N# 	QɅrE*�kVQ3M̤s�A�j��HsD��IC4�6xb�3�A}T�`�fO"�N����F�n�U�p��斃��H&h0��;
��<G$���5;�23�č�7
�ɼ��kU��y��F������*3،YrΩ0��0��E@+&�Vۆ��ɂ	�ĴTZ��32wv�ѲW�]t'&עx��̉�b`w��C`�p&���d)	4�D�j�n8�9l�T&[e7���D��=��%'XN� ��hRf�^eY%Ǟ��{wGUU+�Q?�ے�/�wDhL ��u-��	 �p����#�yIrt*!q7XߦJx�"���T�( Y�����/$�
�1���?�c�"�9
YY�VK8�xpi�ɶT�B���)d�Q�-U�Ổ3��~�����BX���!猜�{Z�VT9���ѳ�~��po�^U��OwG��^�#�  �䅺y�_T��(��̑�r6�	B�Q!%�dk��f����u��W��s�YS��Y�3��[/6��Q��"}W���G#y�g?3ܼ�_��߿0r�w&�%�z�/���^����o{G��cכS�>�jJ�> LsG6I�yD�q"��J�} [  _tc�0w9�\']��9B�DHt�ف{�.k8O
�#�$�$�����] �ٲ���M�?� Ě�ݕ܌:�	�z�P�t�v1�aQL{F�ܤ��~���9S�W0�\U�8qq���. ��� n��+7ew'rnĮV;�ʈ�027�I�9� ��X��lv��~���f^���5��D���>H�>r/�WNNH�N`�5n֐#j�v���LD�w*�+rSm�Zkֱ�n��&���	d�bV-�h��Z/3���݋�X�HD�� D]���̹�W�݃����:w��9�����Lp��^�A�A���;�ɉظ /Vբi�kp�`���(ʒ�����'DH)���w�O��-KϚY�T{�a��B�{Ť`��7L�,+�:V@1��RiԠ�W��������3��$>"Z'�Ĳ�I\�X,���DTHM��b�0� �ݠ�@�7K�k DG߇nI�j�@D� �z̡��H!J�<'�d�)�Ua�����~�	q_�=�	N�����B���Z���C�ê9���K̣+fU@���'kǮG�1�x���`.���'���\�4f�۶(��yE��e�����N{I�<�������c���!Z�3\��3/`�U����b�:�(�Q���X�3���;��z&vx8�=�y�鄾w���<�l�A�O�#\�*����y ���$�b
 l1r�NA��F��Rm�L3yUQ��r�1��R��*5J�Q��:��SͰ�������H0{K\���8�{�F�L[IiˍX	yf��2���p##�A<� V��=O�hDN� �-�_��TGL��Da���;^�=3sΑ,o�c�=m�9���0� �+Sq'*N?%�s"	3�q6��W�:�[e�FnV�Y�Z݈X�qK���qf�� �������� g�VnV�i�����;@�O��DJLF��ff�e���4�p h����Ǡ�Tw6w�AV w_y�/e�����߯�R(�G���į�8jc��o�-��1FQ/jUOO�W�K:�
+��)P��#�  ���K��o�R�)�$a���$���8���ă԰�yL|��	���j�Q���ĝ~��k>�7VIV*��Cv:ξ�b�\=��,GJN_�J���Y�����R~��{�p?�z���'{�Ҥ=��} ��'="q'�8p��=���B9(���A�z;)=P�$����7O�8�p��u�]�����<����POƷ�i�|��v)��໢~7v#����?>W6�L�&}/~�7'�}�ߚ_��[�ίx��&u�'��nF#v4��0	��]�Φ���6f0�=��� 8��8$Np"U�"�)�m1s���%&f%|�@���u��P�fp�LN�`��Y��j}�J Nŗ�j��Ld)�F�1���C ����t0�N���U@�wJ�ٜ�H�wg7��������{/�2���SQ���c�Y�Y��ưB��Fn&�ΰ��Dȣ��+R?S���/�Xg��8��RQ�nK����v�� C�W�C�ɒ�D�_�ލ݀�����,e��� �z̄�z��������V
�Mv�o0	�lP3�X��٬�f>V���=���|�oR�9H�?^��ޠ�4v�p�$�H�2i�������K��c�ԣ���,�dk��_O�ζ���okHǺ�����{$0N'C[���ܩ�ޞ����>K���pd�]U������I?Y*���[8����pc8�5�F`éF�lc�X@I�!̺�EB���p�;c�� �8���[����o��)N�^�����jvv��o'��v8��g��1"�L���Cĩ۟o33�#S!x2*
���($�̂�I�/����
+��Ɉ( 'b#"��<�*͹���dfK���`��o�ۑBS���(RE��?���BÛ��3p.��y;��2�����j11X�L_�ļ<^�BsK	q���������K?U]�9�<�99�嚭?����Z��В��1I�8YS\����f2�Q1��Tw��k>S�2�/���p������P[�A#�\W��-o31�m_�>N�xP��I��0H��'f����VHn)Kލ�H�~ߓ״����u��	F<��~l��G��u���={�ZR��|vm@��i?�|���jWʓ�����Ǖ�ӈߙ��`���-�bZ?��wZ�����~;��BO�N)A	�!}�ZL����@4�*R�Xd�֣�k&�;K[/c{��!ϧʹ��ǿ����`m�m��a��ʕ+�W^�V���7*������~��`ވD mآ��lPYV��l��T[��ӑ��ia+�F�<$ ĸ$; V�8��t��V�&mf0�š��b��Ӿ'Ho#�S���IA. {o�Q��۝A'�*F��t">Rݖ�G�h���ݱS5`+oĞ�e �� ��0�2�9JTa��&ͶT�Ыi0�3 ��5��2�r/��i���i���v���
�^�0�ș��i
��Q�{�nu���W�_U��O�A�r�A������]�OW0_�n=Ni+�`�S2F�����x<�w������jI>9��k��s�YVR�<�yW=߷ߐb夯�i��)\�|Y���*J�����5J�Z���g]I�v�ώ�[�BBP�U��z�������Pwp3�����nF��ۉ�;�lr'�r��o����T6���T�^���t��֔��M�e����<G$�N��en��];C�4ݛ����+����+���g���:�)��8d�8�J	�2����8�s�����L, J�'�P��86�y?Xi�X��i�{�� �B��p�\��J�C��T�ݏ�5+��I_0 �37���6�,� (�w�lH�� �^a��|٧�  ʺt�&/�E�bf,zG����������~�tr���}߭:���!���'�=Y�>��`�Y-��C}*<���SQǎ���)���>?p����q-�u���>P�}�`�U��)��ʳ=��W�>j���B��o�����K�?�D����K^s~[�~ZS=��~@Ik�����71� ���e"��>�al���5Gj����9��(&{��F}��z�0Q4a�?G�b���b,:C��j���4�݄�37:fN�9�����t�
�9����߬_~�VuYh�}=x���E��!��!'CUai"*?|�#�����:KW|� (iQ,��x9^*C�������'/D0:!�����	� �!��2R��p_M����&gD�BV�$w)`}`�����܏���g�c��<~�t_�-���A�S��>q�w@� !�rF)iO�2  �s�{��4���<곤�Ẳ~���~G�vX�!��r2R@��>`���_�{N���QV�J"Z:嗈����X�����'�>��+���K�Ø���K�����$��9
�!��U\����W�e����8�(]k���9?�R���!�]��T�p�Rut���]�m^4�3��5�זkH咉= ���e�=Z�b���!N+�V��P꾟���r����~8�qQ���\y�`���
bU^|�6P�Te2�q����<n��ξ%�e��կ~o�{��]|��L<�x�̻����zwwk2鴍i˃��5����v0kǮ���y��C�Y�E(�Tn���1�ʭ�C�QCZ�..��X9oO�ZH�z.����|eK�B%����0Z��R�A�q����=v����Y�|r{�vi�<P@~���~?�C:�#��Z���)���{U];F�؏)pG�6x�o5�jJ �|�OӀ��o�߸f\!���������    IDAT�$��8�ϱ��ȼt���z����OS?W�'�z�����'�,��`�����a�~������B�\���lҴ��2K��Wa�H�٥�{<�E�.	��~���#z�=�����pߠ�Rڠ�?h;1���e�%Vp��� F@]�`N0� �1�@�����i��P�I�OM�Z������}n����ި~��3D���_���Nr;��h��^|���^�����k�qp��)c2ق�G���Ї�a�~q��Ѥ�:��䬧�� "䜗~|Gj-#�Vsku���;$��$�p�ĺ:���l5��0۲ݫy����$m'ɓ∤�cqL?-I��>,1���պ��|�uߵ���6�"�Q*N>�m���A�?|�S����m�R�c�5s���g��a��q닝��܁O���엎���|��%�{��u)O�<�8 ��9�C���}���x����֚�g?߶������� 60)�2� ����Pw�W�8��$0`��jBA�'u�C!����p0N���}p��� �!���o��k�(.���H�9����`q�+�Ҵm�'?EY�F"��{�=�p�nE�s��9c�"N
�`\J��}���&���������3��úIeݠ�I�yI�:���y���4Y�'�,>_]��u���دo���?����>z��mI�J�w�X�Dq{ƶ�?���K�i��*!Lq��tuK�?�P����0S��������n��o���ݟ�4��;� G�*���V_W_ކr1�0�DwS=��t��s����"��"h��߿{�֭�ǗO��3Y���ŗ�~���/�Qg��������TY��;Mڶ��8��3�w)Y�w?=���P	'�/M@�O��q��� �Xg"|�����>}R����<�5}��w���d?|�׷w�NN?~�Ԙ�(Ռ>�h��j�<<�'"!,-UU��k4M���QU1�Ǆ&61��
"		���7PI��N}��@(�KAd�H s!��~-�չ�� ������j���֎����*�q�ɖ������9���Έ���_Lo���F�����ة�EWј+{9R�1����·�;<��B�G� "ǖ@Zg�|�<c�ͭ��཯��D�2��F��A�^�}>��Ügu0y�y�{<;��Gy������q���8����X�2Ƈ���@eUA����������R��ޑoq��_�w<۝��
�s+I�ѡ��g���fF�]V���SXv$�% �J �$j��Q�FK׉�����Wz���3>�ן��HmB���l��E
���D��.��ю���9�7[\��\�ݴI���F�._���4[)3�_a���<����T�"�Ï[��V[��*���`K����zp�J�;�ez�#��u)�����I�����bR��O���?��u�����V����������ó�<:
�)k�:�O�>X|Č�nB@UU��
�
&,�8	;��KB}%"\�
�sԁʋ�;̙ �LMܝ��9�,-/s�dG�Nd�rMc��7��c���sAoI꯯���}��yI|sF���6��yֹucS��"�#�c�x�vƷ�`��	��,�'}׮	�_���[ �mH�F��ۃ�����ѭ�؇uC��R�;���;(��2������qz�+eyC%�r�9K�{R��*�|p2��4���a�ϯ��X!|�#ĒŬ�i!5��k���T�-H�8�D�2�1�q�T���"sr'"cH�E���%_1�G0�Y͂U���!��S]J<d'�`���,�D�S�/h�XFk��y�L���� kA!T�b*]�9������,�����`�{/�7���?X�U|�O5>R��+W��Wn�F����	o��z�s;��������l7�L�@���f�$|�
�O��9ͻ}:�eb���b��WV�~�C��*���M�q��I������I7�=m|܁�h�Q߯���x@�>�����r�֑�cfNT�B���	������������q����B�ma!̉E2�nj�Djf�UM-#e����]ۉjY�@�ܞL�D�����*檪�X���bfFo����^�t`u�l)���ݾ�Mj|>�g�,��U%x��@nI+&e��]���i-�+_����5k n�i�GD����_U����2���T[����?�n�w�޾��f��2X#�t�-|x�'a�%�F�jC�MF���� ��{q����sr����r�=��p���"~��?N��iWK���}�����G9�3��w��������n����W����Fy�>���c�d�`:ckk�QS�:ƅHh�� �j�9+���������fN9!���Y6�dj9gqgu3/Q�啟lC�Pa�����2sF���AU�,B�N}ri���,��,=]V"��Ւ?\��m����zOЬU�d�� u�!�6g��Q����^y�[���ؘy?�x���+W����V��ua2B�������t���������9	�W�_>��sFJ	A�N��t,��1��P��J2cC?8�01�oOg�|���'}ܳ�I�78����5|^X>
�>��ݫ}Gc�t�U"oG���4�$	�� �W735SS�;����)�T3g$r,�mx� c"���%rd��ȍ9���� �  �3S`��Zq��@U��s�4U誶3tI�@�'�a(�C�ə�劉}�V��� ��VҘe#�T�����dg���>4���D�ݽ[��gOqd�&_��_��\�_���1�zȵՠ��ٝ������c��R:��w0�����
�y/��.'8;�* \��J0����|�n��r.�idYY�#3��Z�+H�ݔ�PZλ}��yq5��<i'`}����~;���i�_���i���y�i�uJ��Nj�۾u.�O2�H�^R�ر��"��7l�jL&4�������%p���	��[#fN #��	� _U�7�5= ���vx+ �|DBu�p�1��Y����تCU[j_��4� �Ч���*
��qN9�9�)�kS<�/0o3�ڤ��� 3LE�vƎR�6f�ˎP��XCUP��Cr��A�x8j�w.=�'Jp%��o6�_6��N�C`o~������3��������"vQI�y�/՘����蕶;����V{0����)��� ���fĩC�������u�瞿�K�.a:�b6�������w�.�Z����~zr���,89��~^]x���6���bu��~�U���fAU���5B]�V71��SA�ٲiVPb�d$���C�]��D��s�w��]�n�����s�������� �v�����?���k�x�G�ɔȦ��9���5@� "����R6�='!"&�:�ZוrS��Lc'�!d��?9 �e�P��8�7�, ��5L�բ�	b�ȠI�"�L�*3`���܅�����)<i��_�����6�9F��ط���]��^�ŝ�Xg��1?����K��]Y�k�,=���Tu�[Q���f���~�~/�������������],�8Β4:֮U�)y4���rR���n��''�#�{i3- ,�QSa<��:��d���]���)�Y��V�_w)�����_(�w�!����Y��?���iFYj���Kӗ���3��a�ۉ~�7S�������}��H��=m�N��*[�:����/��9���McbrS07ĸ��dA���-;)H��'�]�$V�;�Go�-���(��()窊�0������bz݉G��ҿ:����'I��K_�&u�c;a1�)�4�2��^�D/���7ݻ��.u]/#tO��V�݃�y��䏙��(I�U=ťK���W�u���..=?��d
!�Çڡ]d�ԏ��A�;��s� ��i��6�pޜ�R9!@�4>]�=�ow��g>z�x֯o���#j�'O��a�op��� *)�����4�WU�	�"��H��J�� 㞃�5���?���)�Jh��q���X/|��<�ߞ�m��u���g:�N�ƍ�����ڵk����T���!u8�����O��>�į0���>�S�m�6����B�,�w&�ö����:�_hZ	�x�~_�	�}(L�M�$��PW�Uu%�źr�W]����ՐfѶ�	��≑�˗/ǪJ�h�O����\�ؾ���Wg�����/�j#��k�e Ūo��7�i�w	N@
�x�X&P�����jR��C�w�{��-��a� [��4����ն~�m>9	��g�7,�4�PUT̌�|��_�w�>�89�G�_y�+/s��59��s"����:'�@|/�����2�7�����\U�J����W! \U6��Ӆ� pJ[���<���oܸ�� �7�x�oݺE�/_�7�dŽ�_�v́��ۋ�sU�D���������_��k��M^��?�.χ�_c�_�L}������Ȗ���XJ2?,��@��F�����S�V�gAq�����8U�(ֱ�+a���+�w�t�]0���+���� �T�z�ˣ�횦��4����(��������ˇ��/T�
A"rJМ� �Ӄ4��qe�|�f�%|�N�!�1�z���Ӌ�nM����* �	)`1���|��v=�u ��x$��9�V��y�� ���OK�1(|��[[[����|9�e�σ��qj|܁Ow �:�W�{ځROkۿ���x�OWD"��H0OP�U�U�@�ݡ����3�����ڬ`����������ٍ~��^��R]�	���,�(�5��trX����4�F|�+_�����o����bs����{W._�������ƍ �/_0q]���_��=UM/���sq�"�����O�v5���:�QMG]ʵ�s���3sf"g@f
�$>��a �%�,$%P��!"�5ƓI[ג��S�uf�����J4����������-�%<�w�ʕ�4V��Ӧ��RK���-�����K9�q]���03��s03�FJ���3�z�7�)A���8ߠ˜a� � j"�"�d%<w�yT�B�D����A8!�C���T;ޣ���?���u���?����^�F�P���mۢm��ҏ*��Ӟ�?��i�_���9�����������=����5r���*�'%8+1w!63�|Й�:�/�eN򝪵?�������/��k4�ϫ�~������b�@�Q�9���Q��㺙T�d�ĉ��gf���Z4�{��s�����ޞ���/_��/��������������/��a�ʡ5�f�R7�@{ �CgPG����+�Bdf��vPSD$
��㣌�Ď�$]@VI ��q��*����HB ��kSp�Y��W^��t6��͛77��3�'B�&�I|^���V]�"��|v��pߩ뚘�Ѷ-��1��l6�0�L��\q��Wp^ҧp' �5�"����h�!����q�x$ :�3��[3��6<K���i���>�n5��d4���z����������=���=�'�t<����񒾓/t@I�B@�IH�,1	s���~� ���?0�n��>�����ʅш�����l63`��u-�k"��@3��0�ɸ�Z�!��
&NW"�$�:�h�9�d2�w�y��|�M�|�2-�L&��/����� �����o;���޾���Q]��� �Ax?V��l�97�5V�� b ��\-2-鼺sN�D� p��8�����V7�k���J�����[��ao{���×�Z,���9>cx��~��~����1}>��_U�WB75-�/�/��@�BN����7y�,9�;�fo�%��̬\j�D���dG��Ü�0#s ��SꯘO�r���#S�&��!d�[�=+��×�����y�gT�R�,�����#��m��}���jl�ꉦ�K���&�1W�8�ZTŐ�\~Y��Q)PM�u S]{����,"n����2&V#��6�r�%��.��]&�]��QTJ�Ή)PWC����nd$��"��su�6xR��c]���\93#Ɯ��,K�?[�EO�Yz�΅�w1I,Hߢ�岥�v;�:~�+�q�h����<Q~M���Y*ۋ^��B=��̞�}�=���X�w%
�v�����%�v�ųr�˞�����Ҿ����{��O>��%;��by {�����%���E�i�?��?��@K�����-O�QR���H��tx/�W+�+U¨+�ՙ��KE
���_�ݏ�[���t<�:쿴9���ɿ���_������+>��Ѝ|c�@k���S�2UfV�5X4$E!�h`S@C���A�3���,�=��g�{�=��?�g<x�@���x��!�o��?�) K �ө��_���W�������<)�� �w�ӥBLDER�O*t��#!�H�ǻ@̵{�#	o���pf�D�%,u�)\IJ
�����(���r6D��HrZݼ��&�ϤM?�X?��%����X����˕�~8�x���E廱�7ۮ'�.��B& �W���D��D����50-)�cN%S
��_@����ӆ�٬!�D2!%#�\�1Gg	}1ƥ������:�����UbA��[��[rGRۉ�}M��u���ܟ�F�ğu�g���'������/�ٺ�P?�{�>DdA#�iۯ/�^�1��<}�_�<��~��Χ)�2��倫�TQ���pYԃ*y�A(�>�r�D�؝t������D}X9;�"���r��Ϳiy/w��`௪��"U��R����
s��`f1�yT���ټ��ҹ��UA]��VA��Q5gÿ���2���{v��m>���Nj�ш۷o��۷�ʕ+:��h4���?o��"�,����R�w���'j&�L��BũvmG�h/���q��0lH_��l���)$�/�IA�W�F�4ճA]I=(�:_t��d�KH���\�t4��}��¢w0�Bw�B��l`!�E��2x�y���G~�H�耖���!-R��z�2R3���|�5�7�"ZҴ�vi��ug$b<w��J}s�Χ�Yv� �d�_��"Wy��4MKJ��)�|��_�Ó��Y��I�+/���� �.|��=ksu]RxD�s޷��M����[���ck?�+{����z$�f�SR������ӔJBU�eт�"&�m��Sl�R�M:��������������ߗ�÷������EU)�g�B�`�y�y�=tg�}=9�& ��]�����דɤ�'':�yY��ʪtq�EIm���w�N܉+$,qJ�̈́�KOȨbNI_|�RL��������*� �lg�}���}�/�B���:��0��"�(�T`H��,&qy���f�	y��b���8j�D��'�����{w?e0t�*��`c{D]�ܸ�&�yG�%��I��LL�I$�qX&{�Ƚ�ҩ����fvj�[�vAϓ�K\��F�k�?�\�������W������8_cvA�ʲ�����w"�9W�!Y0ѓ$|<����%~��do8�ι�?��4��I�O.�$e�K�Ue�4�YJqn1��Kݏ�ſ,����4����O�@x�w�w���n������M&p��������4�`�B��/��q��b[&�J��ŅXk3���tFJm��U�ˀ�����L=�o���}�YP�d���P%�����v�Νˇ��B���@uh�%+���>S��0�I�R�\����_�{WLs�Lb���`�i���wLg�|����XU��
W����u�̛�d�2o~�����
e1rZxmlp: �w��y�ނ�-��2��]`Q��-�2������l8��л�W�����$K��ئ��EMQID;�4$$$�6L�毛��/���;W�p6Ҵ2��h�r�i ݊�t��u�d��*T]���.���nA������� ����ߓ��=K>��]93��F�k�ʂ(�֩�#1)}�����fBe!�Z����D/�-�������ԏ���	d��B��묒��=    IDATj
�����%~o�"H�Tf� �@x���8������'��'w�G\~}/�mrܽh�E eل����!%v�fT�x���Y_��S�V
VV7�q3qp8�`�������]��Uw�#��	~� ,�<_t/[/.�Ó��M�|ON�l���}A���,}����x�{����eq߽�e��"��!."�d�����>�7�_:;�����:�IUuiY�~�e���(��Ƶ����n��E�я`��+{�'L���hu�b���9��]<��M�Mև�+���z=F��;�R]U�h4�)��e�Y��S�ŔT�,�ixt�\�Ϟ[13�>h�""`q^J<��[���x1�]�:D�h�>�-O��,}O�$�����D�.�jUI6�R
�����1�W���HUU�llq�֫<x𐽃�>RՈ]`y@�&R��ћ���� �ǉ������$8�:�����*�|����-}$�����,Q�9)�Fq>����ʹ���tP��u-�9��,'[U��%1��AV'���7:޹����v�������;X-�0����ae��}_���Ͻğ�����m�d+��j6�B5/g�]ȁݽw�=v�x��]H����0��RBP3K*�daݻ|��x��'`s睈8�d�X�3�>�����$!�"��\GY@�L�{��~�)��̍y����u��+����d82�#�M{�."|˯ǥ'9M)���ey�����%~��h.�b�u=�^3�)����R��y�m��]���ڞ����i~ûr�T���Ih���������	�N]�-��Ģ(���l��?���pؑ>��7�~��"�9�J�5x'V�SAI�"��;���v^���B���B����bT�G_I�\��/$e˛7w*_��\�uD^�m�>�M�'�$�47���I��`�9Y�x�;pa2?M9!��֧QE���"�*9�`��%���
�j�`8,&�M3crrL�-�tc])\AQ��m����nҋ�$����h/��-o�eqQ�/���c.�^��E�]��,iXvO^�%|Z_[>��sXN*������'eٲs�<����{s���y�e�ڦ_7����Г��Y������N�~�۩#�<���+��K�Խ����}R�vP��	�!bw$���l��]4x'�t큨�aR
W���b{o8l���w�?�����-�?��]�r%m\ۈι���w��^��~P��4�:�𾬮�q�bW�a*"&��oڎ�sڕ�
�����{"���
�AL�}E4�dB4c4�`XNU˪t&�"El�0��7ҹ�����r���ⅸw���
��c�0Srֻ���/�v[�&:���>tP(ԑĐZT<b��N9<إ���R�c��7�׹r�%f�#�r|�K��B>�CBw:q���m�8Q�yvY�.��N�[J�4�vY+vѤ��-_���C_��t_�-�c�"�:X�D�@41|մ)>��O��^Ǽ��8�bU%G�,��jw����oۯ����^ 1ѽ������y`S������λ�
����QxM�sVz��� G�Fy4��4M����)K�)�H��,��Kf��@;�L��%�h�b4}�w�ŋ��L�,��">�[�I�����J�)���)��=�D��S���L��y�����G�mlqu{���m,�f���N�ɹ���.�}�O"/�-���r$��g��2ֈ��w>P���w�|�c>+.J��~Z����/p�2��%ΐD��X���d�]A�Pj�k�4�s1��hP=����]�[Yv�FGP�JU%��`.��Kkc��������o	_ j� X
�6��G�?U�êPV�P͊b:oO=O�պC��9�>y{��yz���!D��d2�L����j�r�r��"X���P��h��1�S�p��]|��|�JD=Ε�#E!�4�f����'���������{|���?�'����ō7�y�:u]�
f����O%ςǹD/
t�Ȣ�8·��������$�����R�|U��ǹ���:^���%�E����Z�5N���T}0\4��G�(E��$wp�uM�s�jʔbi�v�4���_����H��B���h2(��{T��)�#�bJI��[Y��**�f�)W�z���AEL%��=+]�	X�	�������5���g����=qV��ʤ����d�u����a�ڳ��jf�tB��Z��C<%��, )�.��HsT$'�4GJs�'�����U�Xl�������k|��B;�0�6�F����N�9*��`�(=Ɠ4\O��=O��]Tw!����=.j�q�b��|��'E_��T�=g�����]�d�T����Lܤ�⯕�~�CZk��%on�������{��?��Ye�nؾ��_���o[�/�/�#W��;'���ʪ�(�<�R/7gɥ����ޣ3d��q*�T0�f����r���ݻ���e5,j�J�����f_b��~l��p���*�{BLfǄ��5�;�־�˱�F�"1u��M�
�D�3��y�{���}�\Y�� "�F#����z�*��Cf����J�mp�u�l�Zvc�6ھq~�͜��ҷ����/�z�h:���z�o/r__��t\�M^,����p.�iJ�rb�U-�|!)kG1�4�Y%���龰�?p���h���߯Zw�?����R]��
@<f�qP�n�L�!K����c&���z��㜊�Unv�N��a�I�k��0<7�[��TW�1&�����$���x<��_�֭[E�d2�������5=Yr9�X$u��라9� �, �9>�����GL&ڕ��,����ƍ<������,J~1��H�����:���"��eH�E�E�_&Z�����/Z۷x_�h|�=X��oï��^�(��C�ab9%HNπz�	�D��Ĕ,&u]w��/Z5_�pD�/
k6�7����i|ݸ>
+��mU���B����[)���,��e��v��4������=Yg��91��/�y��L���HU�n��;�\�o ���5]�E��5��1���ƾV�eI�u������ܾ}���888���K���%���:	�D�����J�ZrTՀ��rxx�����'��+���:����F#�s�S��d��e�ȹek߂�<k���n�/�'���i��ߕ��|���1O�fa�\��"��R�w�K,����ɢE_�����M'|>p铨j�-K�$�Ɖ�WW>�����VnnŮ���V��;gj&�E�s�[�
�h�o;�,*�8�w✊����RS*����ߗw�yǿ��;�Qx�?</��
ZO�f�%M�S�^L��Y���U!����^	�0H��#+M�� �Rp�"�W���8�5�l��}dJ�njC���ʛ���K�)7ߒ	Ww����������x�QY�U�æ#T�(Ig�2�Ѯ�3\���-���:��G||?�ze���IG7����u�+N�#�UX��CB�����(��$�|͋6YT�(��&8�)6��QB��9ae4 !�.��Ɣ�*�2��]G�W�$�	)���dXה*��Z�%|YR�
N)�m�41�LH� BhI��f��Afm0��7D�1��x�D�xQ]�]�=B��GB	(�(f���U5�@�em�fm͑bK�[�V`]��(E�h��pP���`�����ONh�Hj]H!2�$���%�0�Zʲ����|�&|m����nѻ{W|o�}=M;��ܻ�y�ߚ����Q�v���� G�bN����<��L�E�'��FD"��E^T��� uG��w�ύh��&��P�[�-d+jjs�V�9��l��ǜ�R����I�eH��hF�Pf��b�!֟B��GBBp�ߵ�v}PB����Ғ!��G�C��1E�A]��<��N��
�\�H\��b�1:�m�B𑤑 "������.�,�GI��Hj$I�CA۶e	>��Dт.��%j�R��@U1͙�N��k�x�b��༼a���J©�Ԑ�0u6�4���F�릙+�L�a��o����{��J��6�\�t?|�*J�K����_����˓�ͦ��n��5�BKW���T�y2T���H1��D�{�-Ɖlau���9�'�6��>tz�ʊI�Z�|��W�ջԑ�������Gw���:��_^Hʖ�$�r�y���V�%��$�rF۹��Ia���R캆v�B`8T�j��W^e}m1��>��#&�-P4E����B�����4���ܿw��W�P;�Kc0������&m�f�'yB{��X��-/�c��J�B�������Q�pP�:�4����l�t2�x:cg�hF	\]Ǥ4M��guu���5��֩
�w��}�����g�]���.$�]������L�)"1�$e�Or�*/ζwV���b��9�$W����v���u}����eX�z��8:�Ӷ0���!����9�`�>�~�!~�v�?@D�q����ҮO ngD]EP[��G���;l���rf�,�>#������qQ�_tϟ���CDR�$���b��0�$ 2q��dFgж-��E�c� ER��cR���dK��"��9M�[pYV�1&F�F�Gj(j$�#.�G �tr�^�!��������m���yҢ���_�����'�X(Y�H��9�-�B�RD5"^Q�UE�HRC\n�$	R��8<"�� �)R���S
W���fGQ�"���=J)1�:,����:O��̗5���Ec��gfQ̢z�$1o�pH�vʣ*s�L�=t?����}a'���!��M�lX�8�9y�R��=[s�%<�<�,�$b����s"�D�j�hf)��߿.�o��{��?������GL��������eaQF���=v�>U�r)3�'�$�+�	0��d2���{�ܿ��X_�Yٹ�p���gv�p|<e2��"u]0K1[eW�z�	�D� "�63�����2�W���*+�5�_����[L�S���l9Gz���T,��\UYor��67�X�\�\gme��.k 1��89:���]>��3�|�9�Ʉ�:,��Jԕ���1�p��k���k�z�ò�,�{ۗ�h��+�)���@�6��������������w�����w��	�,���O�(��V�^L��Kp����-����[ߺ�͗6Y]U,uЖ�d:�<��Ǭ���o����xX�K'�����9���h�"ބz�M����H�^�Ef�D���8=	����蟉�2AL=�9�0�����:�D�[E���\Љ��D/ƗɞWn	���l���?��	ƫ�|��
������&���J�D��t��p�Zb�������r*�̄����5������e�C�D4!�e�-9�f�)[��`���Y-%0��zo�|!����f*�rZ&�����4�u��Ήa* ��G��>�g/�W���p���DOz�]�L1��s��O���m�SB8ˉ��@"�U]`�ֻe߳����8�""�Du&��P��+dg>E�೎/���ƻ��������_�8�MD$���3U��~���X�N�I$��&̒8����Ԉ9�yդ�h2�����:�o�?z��O�n��Ē�9AΖ�_�b՜�(5�I�G���ߣ�;��"tDli��(|�O&G|��8_҄�nMp~���5��<b��>'�S&��m�fWMO��'}Q<N��f)[v��޿�gkk\���K;#�;W_��˯p��}��'��UD����b�]��k�����׾�[o���[��X��RQy�I�*
�ʓB�l�p���hQrr<a:��R���Q��Q�%W��������;�e{c�A�
ɒm���J�D��хDg�:������m�{�3>�U��;w�����s�e��E�w�U*��>U��A��p�[7_�;����z�����)6İJU�����.
?�iM���g<Nܺ�&��X[����s>��
'�m�	�*N ��}A�	�ق�-89�֩����I�)���]�w6񞒼Ǻ̗�\�*zRG�\m�@�X�/�u�ؿgbɤNL!H��M:{�Eu�t}�29���"!�P'x)p^Q�ݜ�v����]����M|?��߱�6_�إ����1g�i�3�xvOK�{9�5d]G" >���؞�W�!����Tɦ�6Sn�9��Ϸ�'��9���{�$/`�?�GWdKe"��ĮG#�@��|%�-��BL	'�� a��.y�5�O�ED��&��,!Qi���Hw�n��YbE��1�����:�Ǣ�vU�C�}pN������2@_����Bԩ�:ˉ���W�G���.�|�0�K�EM��>g3�#Q����$�ߥŔ�����8=���σ!�pb4�)w�|B�ɢ(����aUS�6ؾ�
/�v�|�§qxrHA�a[�i4��EOnP�	��|:a����L�W�յ-��t���)�=d�Ͳ�/٩��qH)���S��<U�,K���x�����w�ŭ��3('���$u���']���������](IB�y��5������׹v�5���Qj�e�DBgFH�������kEQ��oP���ؠ��/����R�k�Ǔ-��5����^ӂ�H�=�p��K��\���t�	�k�h�������6��P-UA:
/x�Yۺ�`4�HI���=�yC"���;�uH!���N?�O�-2�ҩ<�{.+٪y���Gc���v��[-��M�������!�d�����uvCg��ٓ,��P�:��@�ԏ1[�]�O�ʧ&QA{k�j&��소)[������W�=�_\vz�2Ձw�ښR"Z������T��-�Kz�Z"�EW��j-���RB,��e)e�j2�E�1eˍ�C]�J&X�Zx::��� �9!u${H2�Σa�A+h�Ę�EYP��y�h�/�+=E�yAd)�6�4�K�b��H�w2>��-0���߈�L͂!��ⱘ��W�Y-���o���i��&bD$?7jΝe]83�\���4]�Vg�R����{s��z/�S�n�0uw�|c\��x1e�4&�E fk��<��w�pI��+l!8�~�]ly���3I��C������b2f�������JO��-v6j�шՍk�|�!v��m�MNH*$K��\����(��YJ��b��落�����2�`<������5��'Nf�E�.,��E�Lr{g��pu�j��jM#Ncv�i��󖮝�4{w9>>f��h�&뵊Q��($E9b0�`P���D-�fmG;��t%X�F�o�h��y��0ZYa0,����2�]��|���!���]�/9\|��Mx0���b�e�/kB�bN�ݵ����>L�S��GH���56�����Wj�VG���
�+�ll�ě������O~�t:�=>A,�4�-N-����
��ɹ���'�D>�@��h�x�כ�Xv���]Om5���GJ�.�g��D9d8K�9uX�P�M�Z.����s�E�Qu�k˚y����8�p�'���2��|�!e͞�~��k?S�:����ړ��I2���B,I�X���%�1�]��%��^��\~&GÚ��eRo �Q�\ͧ���-s��U=��=U�y���L�9��	M�е-��u�)����*����>k�����*!VV�X[[��+��$��	M;gz��.[lEN�/�Ӭ}Y�����a�H�%K!�4 �˔$�nv�8�pxX��;u�b�*`�K�_�a�["~}�?5�EQJYV� a�N�N4�>��?|x�)N�K���H��۷=쓒&g��Ÿ���a<�l�[rS�Z��K�I�)�)i3��D�J��a�if�ܻ�	X Ԟ�^��+׮1v��q	��f�C����H@�1��h��I!`��"�9��c������\�2��W�X��a�����C��%�S�ڴ7H��d�G�ޣ��̚�q]��1`\WĶ�d:c���}~�{w�ppp������ߧm��Ρ�A���pEEQV��6U�5S��vyp�{�G4�zw�pr�G�Z�j0b��^�z���V�ͭ���C�2�n&�y�|��FL�l_��hD{7�"�	`JB� ���p��>�����    IDAT�����|�*eI=2����ڕm�]������!��*W���`��������1��N^Յ�,��Y6'8�42TD���)U�yr������%F��E�ʙ'HUz헜Z�R���αUQa���"��k�򂤯� �KS��Q�1s��(}EU8W�
Ż�d�')v�d���ު���j�Eژ�UU�����0��c ����5�vJhbꭔ�E�`KOZ�wc��Ĥ9��N��/D���^�[��VB����sTUE]E��8<4��	)�)�(r_Ԓ.u�%k�o�2���w����l����|�	��1 �0R�'�]��<�������+�5��ܽ��'�E�h8fc�7n������늢�E&�C����}��qpp�H"���/�%W�!j�,�!�R�
# �Q�>~&^�Ǉ� IUI4�L>�"`@]�Rץ��Z#!&	M(�s�{��B1��i[�Yx.�W׵��t�%"9�o������:��{g��lh_�J�'61��B�@�k"Ė���Ķ�XK,
��`m��z����:x���]<���fKR#Y�cy�.��L:,�ل��#hژ����5�zؓ�D�F��vq��u�#n^��:NNN���A�uL�'ܸ����q�����������_���l�rT�s�e���W�!�+�,�e�#�4͌�Ç|����/~�ǟ��d��FO2!t]H���V7���-fM�q�Ǭ�\y���s��O��ϘL���~���ˡ'B�~�(&S�	E&$�&����?�o�����ܶs���yO{��+�U�W�\�Wn����o����:�(hlll0��S5���XZL��w��&�����}x�4��ʗ��_�,t�
KZP�>PDZI�������G�ѣi�k�"!5���Ɩ�����ら�~�>��f���ˬ�����J=P�5E]�R�ifL&�̧��9�����v6��|]�Țؔ���pȵk7x������u�
];ez|���}��a��=��t˜�}!	E֪�Հ��-����rt����=fwwYT�[�Bz�bo&	⠨+VWW������:+�1�~����9��4�H����Sams���|���x��ׯ1��������)���D��'|��'�u�g�9xpb�R���Ң�%h�˯���o��������&�̻@UUl�o�g�����op���S���ݽǝ�?�����l����%s9���pj� Щ���If��c��I���������P\��E�W"-{���A~9�i`�eY�`P�JS�� A�%)���mu���7���e��o������ruSuE,�I2Ra�Y�{1�	�����V��}.D� �]?�)�T��Cb_%aq�G��	]B�H$�w$1b�'���=>��R�z�7^c}|���d��u^y�u������4�)�ù�^����;ʅ�.JW`��	��s%��p��ع������.,�G���<t���eA��u]����;�;����w�bu�fex��h:���G1�Lr����X�R4[L4".��������T>���~�7��_��g��bT4���E�1A�2k#�.��p���m��/��@�������6e�畓�%C�z��/�<a���E BE�T���b8K�4�l�U�"t�޷��<� �I@H���!U5�ƭ[4m��kTU}Z?x:� �SV�m�z�TՀ��b42��ٺ��;9��,�I1�5-��CN���6R����1u=d8Z���fY]]�I�C�����u���(KO]ק�O�L�\��V�ϧt�c�������9:�2�wT��s�S/��W7����3^Y����6k�EAQUT��tQb����{����������î��ҧ{	8�qEE�����o�������IUK��h���}����w�����#U`���D|r���Y�R�cF+�������}���u>��~�ӿ㓓�e���^K�������tμm�Z�d��	�x������笭���l�K&�����pER-!� _���ş���?���q��k+���ks��<m2�YIkc��dkm�O~3��_���kW��!�9�lmo�}�*߽�=��G��@�[7o��+o�֛�amm����ϧ$K�c���Nloƽ{�N����B��������kO4V��;��73�RR����peݚ;��O�#N��$���"2J$ĬO1d��sc�Rt�-��>P�(�Sw$VV%1F��EYX5���j!]�X��R�?wItu�&���[�_'���omŭ�s1r,$�&/�b�­)�q�.+�-m�xߧ49WbLU)ʬ�S���LC�!D�)�n���]�ݽ�����J�)c�\��ε�q���w������k��EB��}^��m98�P��A�+��U9���������a��:����	����f�>�ri� X�t��]/\��f'�A��d�1ϑ�d+'��&�Z2��f8'�pr2���8Ga�� ��8�ݯf����b�{�hh(���Y��3(+�Fe�ꜘ:��J������c2mh�H4��թ�T]q�7��M@�*����֭[\�v���uU}J@;�m|�O��g�?|�g���?c�y��!Z��$aD�V��4������6���:o��W�]cu<ƕIF��S�8��8�EQK̛Yւ����|���_�ɤ��<�/36Gk���k���M�������M����w�:e��x}���Y������ۇ�g�~�����LF�x���Y]]gck���+�olc�cPy��ʠbmu���;|���3�?�Pl�p�hA=�}�*W�^ge}L�"&�ٝ;4M�l�҂�(]�D��`D#�a.��������7YPU>����8�/*:�62�޹���w����׮]a4�4G)�FN=Ml��A<�H�x_CK��-��1{{{Lf-]�9Q��(����D5!�`gg��������_ccm��x��`p��s��Bb6k������=<x�l6���RP��=B���9<�=�>I�)Q3Įn�)�������D����%�8,X���{���B�^��x�$X����������Xx.����8��z3�s�d�l�=z�B�Xʶ�b�E�OK��s[�؄>|��L�'���w5����m6��E�0���]�T5�w�re{�c��Wo��ko�M��p���r`h�R�H�esz��R�tm�d2co����u����YY�dee��f�<�i�����?K�v�09f�	]�S�(r�F\��,��J��>��"@f�,fk\�!��9E��IR������0U���9�MV���˝	����>)j�OA���m$�
�E'BUЀ����� ���,P�!A9j���n��bEYgW�z\�H��h��ԣ1/]���[����os����1������)*_P�R��5�?����
��_����M�����,K�	]H�6ulllp�O�!���?���k�WWr MO2���hq'�z�Eb&{Zd�_j�>8��;�?�Q�
Qq����������z��ׯ�V��AY�Y��5�����@�P�UΏ�uY�N�'��1kZR��S�E���\I��J|5ė�a-lloQ���J�H��u�����mmg��pŀ���y��^��͟���>����R"'=�jf�[;W��wn��[o������~N�3�mnRWbA�r�:߾������W+����4��n��`�(|��y0�:���à�p���������w$s�j�p��xe_V����ޛ,Ir�{~�����1�\��YP @�H^ކ�Lm��`2�B�2Ӫ��3�7��� Z���nKj�� 1՜U��c����8�Y ,Ҭ/�VȪ�ʨH�����N@������p5�V�f:�q9>g>�3[L������S���9:<d>��&	�+N(�p�����^|���/�&(��@Q�����F�sA��������fK�UD��?�m�d�t%:{���xM�<M��tF��s���?O"�v>x�%D|�����*>L��cR�VN��hV1cK�)�=�,��V+�F%,���"6��!K���S�>{-M�;l�;����orvz���*;�#|3~v,��%(DB������t�x��zA�������3jy�?^m��Bo�$��Z΢%�j��뢁��W�|�3K��	��4��� TD���_�Q:�(
�}E���01�!"E�1�g9��+���sͺ��cV����ݨ�B��`��G�C�h�Ӡ�@3&N�,�hM%e]T�QXg��C������;��g��{����W�$x�AI�.��J�f]R�t�nT��NN��0��	(6Z�8�ع�������Oʭ[�h��qL��ZTW�e�"��*�����y�m���ҜCh�r666����w�{�t;�L'E9ie�d�@����0��&K���cgw������\�ˁjQp|z���S���n>���bI��	���k�7TQb�H]+F�9/�/xyrI�u�i������f|9����$1	N��l�D�w��sc��wﰾ��N.��x��K�|���d�B������~�.?�����Z#�R��1GϞr���ň�d�
�BJ�N��dlo�����v6�v��Zo"����fT�RV�����m����~v��z�Y��G����.·L���sF��XE��u��h⬢��O��6]>x-!hq.!H&>t�"7e9��*F?��]�e��e�Y+"b�^y��Kſ���8�Hh솔x	`*�&I^�ܿ��q|�굚�>@AD�	Nh8z�b�����"?��	��&x�m2��5n�챾��.�39=?c>�7#�f�1�V�4����G]MPi�+�<���`���M��6F��m�`��.k�,�b��"7M$��Jc���j泂�tJU
�Q^����������������;�5b�	H�����"c_Or�з�(^V�[E����AB�QT��]���a��G<7(�����a�U;*�s \5�A��A_wQ[5{+�«|��	�ST�F���o+TH1>ڸ�(�A!J�Zy�]���/�.D/�X_�tk�y�������O�m��tp�1��#+���<��ՖD<y�IT���]2��B�E���Ԉ(�����M�~�m~��coo�$m�<,���((˘kt�2:v.`m�s��� �=E9���)O�1�W�J�N����m~����p���<�[Ǽ�y����/�/Jfe�d:��6������:[k=�ַ��V֎���E��
���C|������s��m޸u��A�4Mpa�kT�:��ʯ���WY�$�*���������F> Q���7�����gO(�K��x�#-��������oqcg�V�x...��g_���Cfe�$)e��������wٺ�K�Ip����#>��#?���b�eP��E�v�s{A7ﰵ> ��d-���-�V�Ӌ�_L�$E'm���JR�����ذ-�~������x����,��]��ua��F�%\����~���+|P��H�}Ȕ�\�M�����^zý����s�1~s�ר�\PF<�;'�YQ>i��פ<
(�F7�R���9�	���^_��TP�뵚�?$��/!(V)�MW�'�RE��d���$��u����޽�9ؿ�5�lcΚ,ϥ���J�"�6�F�z�I4�\^����s�n��9�y��.�7vٽ��d6���"*� �K��=7��F�9�x�f��|��)K��G�}fV��W�=V��`S|��-1.N9נs��)�N^N��h��􂁠�C�i�+4����o!�����S�h�5`b�%����EX]^"�P��B�Oy�Z2
\G����H�!&�xoѾ��̅U��M�A��R�G�ΗjL"�VT����=���n߹�;����?a{g�f�(8?�����dBQU�pɀDJ-%��Zl���S:���5(ɘL+T��%�"ow�qc���Gܻw�[wn�j�(���s�<y³g�h�q�S���c�FJ���0"ת�*g\^�svvJQ�h��TB��r��]�}�]���0F���>~ʃGOx��)�Y��(~Q�!�s>�����ҷ�e}='5�4'��D��z���r6gV��rR��]ƣ)�6t;��[x7����ٯp������QB*��$����鈧O�s��.���5�7n�`gs��ጲ��������g��-�N��Y�1Ϗ^���3Ƴ)"-L�Q����6���(C�e�ł�|�pt�x<��/�֓jSq��͠$E�%	"qj��t�����$AJ�$ }v\U�责���9Ϟ<�7��/��8?��\�DE�e���_	/�(�ҳO�`��Q�r�$@)&���BK���y�4|���������g�uxSB���T���[׫�;����%oP%���]Mx��y��������՟��o�X�U&��"�mފ���ky�};�@�]
I${�6��=�֝7IjO+����9NN���8�]fs�k\�
� �����.�y������t�~+es{���999�r4k"IT�͸48$�h�؆=���WYYL&��666�ی�l5Z��(B@y�8�wq̫��#K%t�E$o9b��d(�QhІ�5�ML%E�+t�1LC�F�(�p��Z�H���c��X>D���x���T���W��Wk�<{oc�l��iE�j44���Mu#U1��	E����}��N��`ݜ�Ι/�+��N��������7�bgg�0Ox��9�>���!�јEY`��J6i���@;��{ܻ{���8������9��r�r�hz���͍=~�����~���&y�CUU���~�'���/�#?N����^�ٲn-A�E�ź"�D(Eb4i�����ݻw�qc�ԤX[2�y��1���o9?��|8�v�J[�$A����rD��T6���(���;��+vw�9::��!�@e�x�,j�(n�9�n���D|��Y�_���vH��S��-J�>;"o���;wnq�(v�6������sܼ���0�����}�.7n�@)�t:����|��!�ć�R�� �£Y�Y�{T�o����u�EE(�.M��J���.��798�.����k��D�Ơ���^���΋�>��3~�O����e�yZk�jb݂��]D�}�R�%�k���Z�|[�_w�^{���/���������^6�E�w]e�%H��36ت���X�&K�5��^�h��"���weY�,�V糿�_a�V���tU�:���!z25{�׭���"r��-���`+��Ds~~Ni����Ռ3�`�k�3��(899���)7�{��B��g}s�v;�����j���EH�kޛ֚n�e0�n�ɲ
V�󧨝�|�����B�DH3���z帮>Ռ�B]⛍xxu-��T�Z�(�5X,�ɳ�,K�=�wx�_�����4�n���:_�[>���+�}�k4�$IP!E� ���eFŪ��"tZѤygg���I�YLLg��`��veZnܸ��FDe�G#NNN��ˇ|�駼<:�(
M㥄D�[T��7�����I�#������ޣ�������u�oq�����s���!_|����o9>>FI�l6��Dl���k�)� ����(M��F���^o����v�I���(T���;��Jst�"���9\dI��������&Y#ִJH�k�.F�h���T��J�e�0�/��x��$�#׎�/� �C�L����#=z�����ۨ��	,��^�h��H I2n޼������Q�G�<?<�ɓ'�F#�fZ�(W!:'5i<�"d�6���vsnݺ�Z��%T;��THL�H����kl�]P��H��,Kʲ�A�a�>�G������?棏>�W��Z�h�$*6˸FTuu�,�����]nb���J]�}��u��\KgfM�j������?���~���l�,���[�[7��eL�s�y��^[k��R1Z��t����c�EI\�B��q��R������_|o����z���������tT��G��d    IDAT@�I|���U}�y<�D(M��d�+$�A�����{�TSy�A���Kϋa�f�v�O��ؿ݂`p��#&�)B Q.�?��P�p��ʕx*��0ڒ�0yn8��2�z�<퓦��1;���'�Fl��Ȥ�� m@��.���8&P1] Ҧ.=n1`~vJ���*����7�7�}��W�4�8yV�! ��X�9�c��5�h敥P�"i3��VL�/E�	5$���zM A����$x3��'̫�m��.yk�v��1��$9b��9���.�g]t�&iwy��>?xs�SB&T��8�dt�sbk��Z}���]�-y�|�� ���)Y_vY�gԕèA2D���y}�!z��,���1��8���}�;�w�ug@^ըI�0�����?>���(�i�&�A޿C�o3�Πq�����f ��{9�BSzK��RL`kA��|���޾s��~�j���x�%-��Zz���_�	�������cfG��я��Q��U�����W�@�v !���s�Jpd��&twY�%-�T����������wz�䴶Zm�4�5&�X[[�;H�zG�JQ�9N��.u�#oH�-.��O���EB�:�qA�w0e����N�Q!�,>�H�ٿR;��P8�(��C�R-9E�K�82���n�c��/����_�O��O�͵�}�m�j��=Ϟ>�w�����o�霾�(U�I�p
�n�kn�z�����,ׄv�{Xզv��VD�Eb���yYF��Ω�0�O)JC�Y=��s��>�!e��nVq���|��#g���}����3pe�$!*�E"��-��K���ٔ)UƽbPT.�i�`�ޢʂ��V�٤���R���myO��>�M6�zk4�%�0J����x����$�������� !�R_-P�N���D7ݸ`�f2�V��I�N�T��i����4�*����� U��{��T�uJ�%(�q�k߿��������^W���$+h����9��e��O���t�pt�h|�V�&1	��W3���G�e�t6n��$�¶���D��2�]`�������s���m�ӡ���v�S��q�k
~����*&�	��^n�TV����Q��^�}W���6O!�t��F�h��"o�ź&p]��,gms��7�*��P������Y	*�;�`��>o������Z	�.�8;�уǜ��,\�����ӝ���r��E���������{�E�t2a:�b��V����N��Fb2��n�fkg���-�<��/>��,�9���DY��Zk>��i���W�]�VƬ��,� hu2���mm���esm�^/��G��GF�	T�bQ-�\����ǰ����������y����B'h�%x��ټij��ڤ�A$���N�,	�vމ\HJL3FLp��IIL���Q%"c��Xg��1q&X��K�窕�,ƀ�
������چR�w��MC|��m�}�Ngc���8�ء�f�6�޽���g'����޽��۷����9���<�����,3D��K���@�V*���	�3�qd49�$��qA���yJ��Z�V�6B��|��%'''��q)�h�]���0�8::����1���V*+����{��4Z�$�։�i���A1��c��p�>��? >\������'y]�����n���@��R]�	ޛW����4��5;�oqz�#z�d��6P"�9+���?��?������������z�����3���6!��	���Ңoy �dCp� �<�W�'�����숃�,���2�Q�)����%��S-ב��E�ƍW)�
,�.	v�h4�����l�n7#�r��y��HL����(_�����������׻��j"ˢ9��5}���w��B|��k�RB�bk"�|=.*,sa�HX5�}�E��e(T��������`0��>�$�h�|^0��=�[�tY�3N�^������׿��0�s-�$y��t��W�p����4N��K�B`<q||L9_0�ssw��`��"{�>y���pȳg_������?���xF�b�%(�,���'�s�v�fk�O���LB��1��'hI1�Kj$�Ҿd^�Iۊ�{�p$1^,$i	�|���QQv�iuԊ?i��:��<ĦPC��$���h�)Y��q�uAK�vY`�����Zu�u��^�H�;��c��Z.�%''_<cVN����j�Ij���I�ZX7���ԾB%�nhiH&1�f�p.�DΝw5"	���
.��8|򄃭���5�z=v�n���?"Ks�o޻���-��.�ل�O����CF�<Y�!1�9*a%f��`�!���5\ښ��S,&T�ʥX��ϑ���xo�
噌/9:~��'O8|�yQ�t�h)-��4���j�q�"�R�R�D�\������%�����u�*��	^��D�J�ȮJÖ��y�ˤ����{z���/~��W����?���h<>Ͳl]'��^!��#ڈ��Z�e�Ue)W}KaLs���t���M�r��~��1A+%Ai��!�F��y"a������TR��u͙������IxM�
�L��S���b@y�R��huKUL�O9?;b:�E�B+�HҢ��dk{���\�_4Q4�@�W�I�o0~�1pVJ!A��QU%�٘�x��fT>.5��.�:�+b��9�@Y����7�����Ѷ�Ղ��A}Q�xƇ_��ӫfԣ�Ҝ:D�x��(E����(e�Q:�3X�~���]�I	�Py!1-*;DDa�6MB�縺b:�ɯ������3f��		����_v��I�1QMmd*D�V�E��A)E�=�E���;;[�Y4^���(�Ŕ'�>��ɣ�py�t/��/:`�x(}�����,�2	)�)tPh��i�D�_'�x^N��iQ2��)�%$����c�b�Qe�!(�.T��:�o�77����`Xb@�53�f�Dى�%&r�$P�|(�PTT�)ò��:z����U�s��ZB������ٳ'�������!H�&�A)A)�ҁ@���2~t�6��B䲪&�'���ޡ�4"�D�S#xWq9<�<}��v�[Z�6��?��w��更RE����b��/x��g�'8_�[,:�x/,=���F録X0:�����O�YR��-XrjU������+�j����t���H�I�ީ�z��cV�E]a�IB]�WԐk�kR�^����υ Uei�rc�$A$/-A��}���L�<TU!�^O��n����A���T��dY'�z��ӿ�ȏ�u��%�:S�eVV���9|Ղ���WH�7Mv�
lcB�""��
<����+k��V\��9��#>D�Y\c�-#iUK�7�݈`�EU$�;�lz���s��ȩm�h�!o����e}�����$����z����2���_�o=x�r�p8d:��� cZY�~-�"B�jJ^ݑ}��s�f��`���L��n��x3/�?p̖���j�7:�t���л�T� �HZ5i\�y�j��q$�$	:i��Qdy�v�M���jaV�(�Ap$IF���:PU5*8�/Ny��3~������)�t�Q	�����I�&��x���hcل(Qe"�Iw)��bX�ɑ��W�`H�൥���Gǃ�e<<"O*
���:��FH�xm�����<Ƥey�Ea)m�V��m��*�(�0Z#�B�cr9���/N^2�Ϩ�8*&Մ��2:4�Fŉ!����
���� <4~E�6�RsM�(��@��D�T@+��btq���Ng#��Z���sM+���|�t:���X׎����.�gq�e""�Q�DB�Fi�I&�
:U�<���m�����I@�L�J�&<�q�W�gCN���O;dY4��Z9k[�l-��������/���Ǐ2��"(�ƈ�#^����
���E��<!K�Mk����G����C&�&ic���lؠe	Ҩ��5����(�bm I�>>Ьe��kJ^��*'4������Z��U�A�އ�u��e�
��
��V�8��7?�:yxy�8__�닋Too�rx����;Q�����!�j�8rJ����[�B?�1ʹ�Tu�TUi����s��2h��
��jσ��}���B*Jk��VB�j�oz����^��Õ[� ދ���-[�W�9ML�pED�DS,.99~�'�0��x7�t����8�h��u��J��l���q�4&����i���l��Y�,[tL M���}�,g6/vD�b�ثuݪ�V�D��׵t�ո:6�ZA�#��}�`�J�-V#��AGT��f�7F�e9�Ic"��h>�tT�zE�^%�i�Uѧn��c�(�1:?�����GϢ��GR!z6�i�1�n���5Ƭ·J���ʢ����GO����$o�u7��v�R�Ep5�ٔ��3F���bM�C�9�I��k�$(�N���삗����<!�:EEQV�N(B75>AH��_I��H�x����_~���h�i8<�S|0(�V�N�G��f:)�6�/�ll��1㎈���(Y��b���hţ���|��ƀ��aK��hƳ�S>z�%�ш�l�B˽�C�A\U�r�{�L&��c:u�%��(<u��h�:�IS�iP~H[1%o{��x[�G�(ݼ���K�; ʡ�`�soy���wYT���$�:�
X�N��t���S��O�m��$��x����@�%�ɬ�U[�<#1m���*t+mI�
	<8���_c&�u�B�����l�٘]�VYnڜ�]կ.�W��oF����~��)x��DEDi�m0�����|��ϊb2�v����)��]z
���� ����4�x<֭��ot�_b+%::ŖE��L��^�#�-���"�z�[���h���XV�l�F�Ң�(Z���������^��+ct��]�Ba��-�4I�}�%M<��-0J�U��&��{F8Y��JS��M�6�������./��!�$��ɑƻ,6A��Ҟ�.���C��Nא�ڬ�Ek��0�̿
��~�k�f_�����ﵓ�G�xdV{s���+�/���j�_q��o�b�4#����)�ݖjN�5&��Яb-�ق�dĢ���5��k������������UE1��'��Z��ʤ�������fιՃX)MՂ�d���3�=����q9��]ۤ�
k���HM 5B�
�!k����`�ńZ"oL�mZ������
cbsrt���G̋���'B��D�^C#
%��L8*.�#�ʣ��Y���xhe	��wnߣ\�9>z���|5&�bJP0���L���a\�XB��傋�S��Oh�����o�L�V{�2�sqq��:��@ek���.P���
-�o�˫H���1'8�b�b�=`k{���]���i��Q����7�X,JNG�J�5�]�������z�x�s�P3��<;z���ǤiJ���h�jŕ����%�|F���q{�F8��F�6F�b��b����t�$�ps���t}.//լ&���;�6�t<f2�dQ�i���-���=K�]fl+uM��$�HC�_�ZYZ.5�_���⻖������	��|���S�|��I��Å�^�?6J��'������f#�pz�~���?��������1���E9wO�q�*+ŢJ�"��f�?���V����^9Y_�u7�Ʒ�9PJ��*4���('���̿���^/��T$	�DB��κ?jIY����Z�W$H��ؼ)#TuE1��=�����z��\#��m�����B�eE$�/я@l�L"�V#���Y�I�����A��g|6�[�v_�.���\��;-2�F�\�7�^V�+���b���D�E�Z,V��Չ�ʸ+�4&�:o�����(�'g'<{���'���1I���6n����{�9I kKL�$&gmm���5���UAY.�E� 6�������r�~}��\�x4���!���>���#�<IQy��;�c�bVVܹu�!K2Zy���Lo����EM�
�3L�ct�w��t�W�,�X__����z���K\ KeI��rV���x����.��%Y�C�d*!x(��ɘb:a1_���Nw���w)���Ֆ�\D�OPH0� ѓ0�wK�P�ӨA�;|1'(�r���/��i�LF������~�ڠ�˗9���6 UUD��tJY,"�aqδ���B+R�!h�7qC����&a���`�?���w�����bm}��o���t(?{@�X0����b��2"�w�v兠^�<�����no���Gy��f��<}�gϞqzz�W+iL��xo���q5*Tԕ0�sv|D'KI�gm�����n��[��ՆO�Q	Jiʲ���'O�����OYT��}�Fk� ��gt�ED_�&����B��Y2z_��yK�Jϑ�D�jU�E)��4�`���Y��cv,�0׋4mϒ3��(Z�V�_tC��{�%�On'm��u���d���Jkkq��lj�Z�(^�̷��~�K�~NW�h_�zq)Q!���Q*�J�|��߿/�����>��C�I](iϕR����ת�-�j!J"�D�х�
ثrt������j���>�B������^��;o��BQY��6��������S�D���$11!�l�Ѝ���c]�u���
7&��h�������6�OO(��t5޽�9Tl,E�>ٲ���ż&�ID�p�nB]�e�FQ7�Ө��RW.B�ί�4�4���\g�'-kG߾łn�����[c2�EkMh�8�[!r�.U`y;糇���������i4���<~��gsn�Ϩ����M�Y���N��O~�3����#·�r��Rʪ��KT�"�߾��![�&f��g�����j���)UU�����������W�LQ:�פY�|1���2^�xy�_Wܺy�V�!o��w~��`���]l��	E�qV��Z^�8���%7����	���m����4>��cF���b<�ɵCD�%Q!�g>�1�Ϩ���ʨm���ʒIF��|��G�����"�Ak���]�Ii�Z�L��s�kOYG��[$IF�g-�
WVL�#./ǔ��	�����c:t;�l��i%}���u�w眃��eI1�9�g5u]3���8���ϟqyYPۈ�4A����
��߿�_������{j��1�� ��ǻ��=�{���7�կ~�d2i���,��6E���,퉪x�7�[G�Փ'O��w�~7��2�jA����?��������@�c��JҨ�vok���G_|�txNU��[?�����N�v7G�h���Z%X�wn����V���c �G���ʹ�Y[�S�\m)˒�dL&��ycU��i9Y5����7ڱ\kJD�r�p8H҄�*�i��I˪hk�Z���5�����>�&�����Lc��A-���i��m�~�ӟw������mv���o���m�H-BR,����$�$"�����<ֹ�O�r��r�B4�.�Y�IL��:��H�D��!��K�����A��������㏿w�(��z��������T.B�^��JI���?�u��fÑ�*�X��=k|�[TH��cU���/�NRҴ�Z��HCr��6�*ߠ�}�_I�Ccyʲ1�C�q_�7�k-��R�S�Yކ�xl�ڴ�4o�e-"v��[]Z�i�am�1M$MS�xW��BՃ�B�f��|�d:b23�M(�cQ�S&�F�3��9�op��>�kk�SC��S�9�]0�g\��P�|�Jd��e�z�*5�?G�j<:���R[����{��6F<�d�~+gmm�v�cm@K�����zLU9jU1�8=>�r�&��6F)��6*l��[���	'g'���,���"�2�&�b2����K����F�}7v;J���3��x���G_0�[���u�t6i�Z�:]n޼I]͗S���#ht-w*q�y(�)Ǉ��򋇼8���<�W�e���×t�5�Ulml��{��ݽRH���*`m��5E1g6��P��Fc�HL	���J`�����wx덷�ٹ� I ��*xt����l@Q�x�����1�$|��M�5/����?3C�    IDAT|Nϼ,�ᐧO���ssg�b>���Grޠ|W��cL��Fm⫨.����kz����~/GT�(A��zO�bڈ�)�^�;N���H���+[��<*(���Ղ�t�h8$	�Ʉ�(V����=4��_�{�[}�9ޞ�m�(z�H�E�:WՠL��R�?-�������ԡ���N�]�>F���_\Cr���W�ͺ��I�2���j�V�.�^��)�t>����|Y�}=��g�sN���!��c��ޙN�-����Q�V�7�L$s�
�t$!.N7��*s�ܽ:�kIĂ�Z��o�# ����j]W3��V��@i�E�м�u�Ĳ�[�dF���I�������[��{Z5�ߡ\"��g.���G����vz��t:=�2XOK�u�.��-0]p92�Wxp!�s���F���h�2��m��(3\]���Qc뀳0�O(&c��PԴ����f���O���NY�������PB���},����$^�Sj��[��hmQ8_���Y�!��;�yA�:X�F�w�X����[@r��X�̊9��/.y��1k�d�a{��w3L����6;��<9|F���5���V��D4x6���S~�ϖ��W�	*$�ה��U��&��D��cs�M;���ln�@�a�\|�/G�"8-�U��P-x<�3�L8�Q5�ʨl��r�cP�������Q{{�dgR7�  8D*���m��6�8����J�A��"��i]�L��)�����;�i����zl7mJI�C�Ao�v��{�#%(cb���jWOh�J������|N��{����?��'0	�c����L"��9�&x��������g|�EME�7����u�t�,n]���b��H���999c8���
.
��5���������+馚Ǐs9R�q�-J}M+4^�&�Z!P�:ˀs%!h���u%J%�uκP�Y�1E�MI����i˟�I=i-.��M��+���?��%�������� -R�VR�O*�[��&I0FW�z]����t��u܈E:�%Ѳ)�_˧��oЬx���9P[+�7����%"�ޫ���߿>��ÿ���[��W���E!�Vˇ��b��I{���X��~�<���k-�%��ɞA��h�8tX����$�J0є��W��#������o���1�
)�}u�DZ7���t^7On�Zln�q��>w�q�{��khӂԢ�܂��\pt��O�����c���]��ǋF���$�	��5�h���e�b4$ʠ�`E�XB5c|�ç�v�`n�ڦ�O�m�r�U��x����!����.OrdYz���{�="2	$�B�����j>�j(3Y%�43iQZHF3��h-�?@f�ϖ�^i%�dM�E�#gĚ~Uw=�F&����p����u�G"�LTݨ�<f�gDFzxx�����|�;8'�Z��y��:�+:���@Dh����.��k"�8�()5�Fxx�KJQ�F��-n�{��[(F��o]��u< �Y��Φܻw���h@�{k.R9a0\gta��I��̳u�*o]����y�i.)K���+b�kc:K�-�R
���p�.E��2k��oq���
�A�\p$.WxӷcK��V\�T%��P�%B64vE�,m��'O1�[��1��1���[����1���ѣ) 8�S�x��)�qC�b��� ii���*�f;����vΚ��T�6�͘��5����_��3��w>�l(�X4�o�\K�r�d�	 N"F[�i���	�4���G����翡��	��5�!�c���QV{�RX	4��wwB�3&�k�qy��!%�@�az8�����i޿˝�>��'�ۨ�
Vrߑf�!���/�~|��Qvw�u~�)W�΋7�n��@]f���y�����2x/�HmLM(lBJo��?j��vY5>5F+�ݵ����O�d�>�� >�����O���G:�����b���+�;�Ժ�lTIM3[�����d��nE��ub!ʏ�Ʌ��҅1�X�R��K�����U����fę@߭���(�h�h��4�XPe���x_�j�[��v	����:hD�JT$!��p.d]�vI�>��ٿ*3�9��e��-�MSVD�$��������2�_ЍkG�
���tU�!d�6�r�*7?��?���~��K��k����^�����m��u��K�؟Ly�7f'9M���p���:��m�>��|;����fF�5��A�jIi��<݆_H��#޻u��Kk�oq��m.]��<��g���K��|��[�M�Svww���c<x���>I��o�BR�U�%�{;�'f��{4�6��������}b�`�$ib|���/͔0�0���֥.\X�	��X���amT��ŷ-�ㆺ�D1�u8[`m�e���0Fi��w�&�;�Ƿ��w�z�2��̩z'�2�qX!j������u���N�o����SNժ�t̠OS<!Lr���{̏��b�!�������*�������|��`>*>v��C��Aei�	�}�k'�lm] Ě�3��g�lS0*���'��<�������,")֮��F�O�9/A�$�~q����}�t����Z�!�-P�`M�B,��<%E4`D�.���1�����1���s�chĄzU��[bPJ��g:�#�Y��I$��ɴ��G�-�l���s������b�S8���Ң�������=Lw��1�oo��n(Ӭ�O�̧G%b�!�j�8Ve]Y#�u5�����4|�-��?�O?���~?����Xo�������9��5��4�se��PO&��'O6�ww�tC�EI����en�u.��E�6`�qh����%�
"b:џ��T�L�1���/������k:5��ƙ@_Bw��H�B��=]~�E����Ӹ�J1�!�V��Iٜ؂+��&EUs�*LgP,���с=Y������������X�SY}��M�:�[����h4����|��G|����z��%$�Qm�M�ea�8b:�Y�ؤ�z���p0�&�U�������Y]���O��6��^��2@�1��#M��$0�3����8�Nx��7ih�7��i�u�8k�i���Jz��m[f�>�W��'������石��Z �^S��)O܉�H�	��=�ٲ�����C�Z&��G�~�d�MJ�%I�D-��{�l:�`o��G��y�W�^Ŕ�<`�����ȓ�S.]�`4rԓ=?���_���~y[s�-�C�%�W�t��<3��9��������;��F%X����Z+m}H���N����.��?$�DU��5��
�;<ԓ�GgL�O�N']Ex���͔�B�ޙDY8o��`o'�EM�F��)����������{��x���6�g�4�Y�+^�Au�?�X�f:�Bw~����Ε,*��\5�ӻ�.c ��ͨ�MTeA�a�k3[ �n�h1��jn��'h�H�"m8Z��s0> ��ԶB4g&��ۯ��x�YM���qHS7<Y�I����b����|��|̅��
/�=+z�X7�	��x��g^�+��j��j��N�)B�FA���$�B�	�������8Wa� }��'|��O_A��W|�O������'�Z;M��ǅ�ֶ�ș�Z[��¬��{{����Ҷ-�ᐶ^tԀ�E2��dڏu���L)�jV�cz.Ѫ�aT.����򓟸�
�oO��FkL/������Ǒ�2a��K�U�K~~�ӑ�ib��e��{�M�����E�tMy�:��X��I˞ږ���o��	>}9@QW� tm���Cd\O�I����0EC��)���eg�)��Ɏ�H��~�ij?~̯~�+�<���o���ϙ�p�|���"b�1B
D��:�������<�~cZv������LC�s�ٳ�,9���f�����p������MӐb���t�Q�&�B�S�*�����=�pv�W�Q&��_��S��Tw]�[���L����s��}.l^"Y�`<e<��g}�2kÒ����gw�.O��gz�K�BU�C!�x(�l;�}�8RPB���f��?�*�)�1������|����~���� _?%�O�O���Q�@�DA\�X!Ɩz6CS��䰻�)6� :E�DDsG�f8c(J�T�^hSM2UK݌��W��!�m���o)6�EI]7�Pж��aN���C��RN���C��b��ռ�p��f#]�UL!��8����:5�K�gP�XbP�5X1(	M>��IH*X7@����b�Q$Ke�0����̅����-޷�~9g�j����]�[�����O���c����is1/��: 5�b�y�W���fw����[�1ѵ6�V�vXɪ��Ŀ[8[��u2����a8����G?����_���'vs�q��?Y�5����?qI�'�A1����4m9>8ܘL&.�,�D@��<�I��Y���`�8�f�����#�N��T%�:��lc*���*$����3���s�U	A��$Uc�(�|��E'�~��S����C6t�Wg.����8�V)�k(V�#���2�޿��8�qٖ��U���~���k��o<��_���t��*�k���f�	|M�cB}H�v�<��d<g�g988 FK1(1����;��1���~������|����6t�-��Ɩ'O�p0>���#O[�3���-W`��6�:�_7��V����>١r�������JLk:��k#�@��hB�p�ϸ�	dm`)�!Ea�}"�-e�!J[�����c\�&ԖH��!Q�1��Q�QڀȄ䧐��I!���1Xk��@���)`�Hg:]O�k���r�)�Hf�А��Y���2�m��bPr��JT!h�$���qW!D�`�v�#崣��H��F���lJHu��i�mZ�R�1B�&Q�HDf��WLYfB�<�u�o�o�{q���,@U�o���b����͆�JW@�L�����lC��l�}�I��M1`�ҕG*�mC@	����{9�|>F��F�9��YK���/:0I�d޶-V���H1��L�;|\��*^���>�;vrn�[D��Q/�$Ĵ�
{�IBJ~�!�XSUv�&L��OJ�X����~b~�㟙���gG�1������V:w�R�ܞ��c���z�Q U���Q�g͠���Y��#y1*2\��qQ�x�X�Or����j�uSծ�KlLq���`/�n���x��,�O�����L�V�q�&��5	�N�-�XTɓ�Ƣ�U$w��<,�Эf��)�m����Z�F��lfk
<-�Xc+�t<�Z�����%�P��w	�RT�v���e���>`K
r�1M>8�*�4�1�3p��{�7f�ʈd*� 53��Sf������}�n����1J���8��!�<��~���se�*1���ȣf�)I)�6?15����ȕ�
�1ⳬ����;�[��bp��J�9Mn�RPtm':i�j��-.�rv>y^U���sʪB"[uV�i�c��l>/H!Rh��~�ՙD$c��su\�P���s�6B؁�C�����>R~}вh��#��0L'm78J�Ďc�1� ��@Y�m�����'H.͏_ �ݙ���EJ����`�J����:��^��t�-�o�!Q0���S����k�':�N׵/1�<g�.���UC*����I�4�'����˔U�82��{D��k�Gl($�^#��WgX�Ou��EP
F4��巏�Pu��q.%%H�R�5�[�H����I6W E�y���\���������7)X�)�|DT�K�f�W�RJk�&R��f���؋&��0���J[��+��O�n�?�ѧf��j�w�����S4w���n���'���R��*�K�1�}%�������U����d�1�r������A�ˆ�>t��������?�Ʈ~iI=Vk1)��)ϯ��Q��L��11)��@���Jj�0Ŗ�%v������gc��U:F�0&%!�u1�d����u�?Z��7�JB��}CU�y���(�������EvN�/?�wqH)Q75�{{f��q�����n�V�����
!t��ɼ[ċb�ZK+������r�끗�*(�"��B�٪Fcw� gW����i�$���V��G���O��8�~��U��*Q�:H�Y�;c�F�����Kg�.�5��O�wf���p��7>�[Ě�K׸������>������I���6�E��m��(T��!������]Cz�0v�XhQUuRu�Y[M7�f6�!�)��d.��^/Y�u������t���y��������^}ߢ8[!�z�=
'�ݚD��d���_�+8�]��Z�I	��]X�8�w�����S�5M�d� ̭WV,Z,I�-W�j��X��+2@��<~����]BH81E�1j��@����!/^dss�A���0�����$3Σ`����O�ǐ-d�h:��B3k��$�:*5��XYM���2�8
0^%�8�����*��i:���y�&��͓�����1W8ۈ��v���%�d�q��GEQ�����ч����_�6������U����pq:������z�O,l<']��'��>dk�謽��dR��ު�쟪�7+����!��)�Z�j�4�l4�N7Ƈ�E�4Y*�V���ŽesW,��E$��I�(DT�ALix���'v^��-�3rlI�HL;/�:s,"9����]��RM�QJY���֗���A��>�X�*@c-�a�h4��+���kvvv8<<̀�Ȃ���t��]ڼ��o��[W/�6Ќ's�O��B_|.�Vy�� ��++)!��*�3�v��\�����A�eA�:(8��������5����?����o��=��~˯;��N0�����4�+��ê*�Y�F�U�O�[8�/[�M�?+Fͧi���TվrՌ~��?��ʁ���w����?���>*q���?�,������U�+_i�FwyjL3S����b+�?J��7��w<�[냑Sgdm0l�1ƇP6���Y]�O��y�^�ڟ�Si�_Ac3Ţi^@�C$��%q8+��ί6���<^y�Iӷ���$�I&�K"&i�����`��;͕&b�nA��� ��a}m@QX��Q9�og��<a{{�}���x)2UE����K��" (Y���>�r���'�������VX �$Yk��9�|ik��׮r�������Ã��2O�+����N��F�����lQ#�pe��>-���E!ar��ף�>�W˓�d�NJ/����4�uX>!�k�$�F�Q��j0��?��sM�j ��i�Q.���p�P����Ц;X�����׳bˇR�n����z�%���vZb\�&4��8w����}W�vW�ߨ��ٌ4���������
6S9*�5�~���v�b�Δ�rMqV\ҤҴͰ���tR�,S�[u���h���~��@5%$t ��@Hڦ�T��^��|����:rxo�Pp	�6%HJ�uH�9ӷ�^~*ɵ�BF0�!"�͌���\���/_b8(�~��Ç�~��z4����6j}��%�b�K������ds�kX'�f-��v��E��5��iU��$B����pĥU��qx����cU�'��42��v���i裐��T����x��_�3�|���q����*Nf�~w��� �o&�������災��qϩ*Ei��i"EQu�z�m�Uj�Z_ۜj�֕E+FRR5)�.!}��	�}��~
��Y��^/�֤Cm�P��G�!<����ڎ��ҍ�{ab�nĢ�k6��B5ҡ	0�n��6v͖���?֔>H�ه�UAGU5�UY�\TM�o�Q;�mx�}�ڦi�v\���(���&^������R�c�6DB�F�[��y�o_�	�ŵ$d+�؈:U5"G�ď퍗{���;��#����"]C��K|��;���[\��"����Gܿw����K��}ȕq1k�b��(��P5(��Xc}4��'���=e�`/[6��y{�{*ٹ�ϻ ��    IDATH��Z�%���鄃�]���2�N�L�T�����Aa��i�Y�TL6}�k��1��'ѐ�0Y�>\���4}��e:���E �U|���y�5^���_�G�"��Ѣ��N�X��DFeYVj��� )�PT�ںn�1�^5����$�=I�`�Rnc���ZQ�E����jU�q:L��D�Vn�GFt+Z�D��tr	�+Q규wkɷ�c���n8W���Z] �@<���:F?�L��I����t:z��|�nKO����{��.lI���FB�4��U�I��1\��~��� �-��i��(`�}�$�dR�6�/T8Q�Ē<��1	���)Pcx��5޻}�wo\g4������#�>}�o)��ި�8�̲)����F��P��������YSO���:#Y��-��N0I��b%kg(��Id��4������H52'}+i�#^ F�bD���J�W�e3ꤽ�����w��v_���y�&��b�{�%215�Y@U(܀�pHJ	��_��E��u���5]S����R�B1�)�!�Ԋ�Z7j̄H� �u4^ ���v]�#����)m�&�a��� �c5O.���cw��/��2��\��-��\���E�����B!M�b�{�F�|��?8g��MqЗ�>.�X^�d6E�PD�pe]W N_��wOP�ڳ��FM�2\[����*�!�W�)x��w������7x��U���޽�l?~ȓ�;��I$�eF,���	[qEE�F4m�(,�{�ׯ18,���|��_�gUU1�L(\E�b!��RG�+��	�ʕ+8������W0�1�\~�׃,�
  ���������r��Q�ٓ�2 㤮"�������<�D�wg�A�	���q����}6�s{���,Kʮ7o۶�I�vZ���/�����糂ھ���kW�ɯ4��L심YN)冚��Wg���.8"٨:!�h�����{ՠ2h�j*�"8gP�2�Xi�/$R���V�zM�Ψ �
�*;�ͫ�%O�����P8�jJ���0�8��l4kf.���s���ׇ������;�eM{	UW���}v�(�K�l&�>��\>)�}0���ӟ&�����[gb�Jk5U���%f	��Iz�>�~�㪪HbH�-iC.�غ|���y�;�x��UF�����}u�P�5�]�_�N��j�blژH�FL�ŋ�q�m޽q�A阌�9�ߧm�DB��ш+���u�(�BdPX��u6FCJ� �L'�L�����1Z��	�t���fiۅ,�Wo��t�LC߲k828<<<����8�}.sx�at1$r�a5��<��E�)x�Z�h��(E�*I��S����El0֥���8��AEDEcD�dj��q��)]D-�4u�&��!�!�*xoC�4�r�Ƌ�u�S�����Q�1j�Qb�x�cw�)��MN^���`�ٲ��ֺR���}A���XN�������!t�Ƹ\�Q�z�&|�޹q���!m[s��W|��_���}f���a�D���*�������n��wo��kW0ֳ�󘇏�3����1FhB^iI���GX_��z�*�/_f}mH�3&��1��H)��p��/��=8�Mq�r��z�
����8~9zV�(���k:�3�Fͼ���~ Ů7�t�|�ShE0�řO��[�5bR�)*�@JEU4�I�Ģ�k�.�;n?+��EPє��dU�A0�{������p�{s��߿��Y?rQe�;���\��N�<ޘ8�{\�+���M!/uu'����5Ε`
\5��[7���l]y��2LǇܻ�_���ܹ�%��!)eX���	\��� SW�+��pĻ�����=�~������{<����l�%kQ��I�jD�ź���$�j�ƥ�Wٺt�����a:�g6��O����g�!���P2�v�v�V�|��Y��x��h5e�c	�'�E�ӋS���X>7G��]�����}�CU�G�f�y�Ҩq��������+FZ�5	�$�FAS���hcD-�I��,7�l2(J��������rG�|���ӂ�ש��x���`�1�<C���!�կ����gf����RKnM�]A�Iz���j��h�(�؂ \X����~�ÿɥ�ˠOy�����_����<y�M���j:���C����9�5��ܾ͋�����ryk��-���<|����'���]���U@=V�`�)sJ��`\6v����>�Oi�Iw#�\XqV���g��i]l�	����c�oE,�{��ih�����ى�П�k��+�����-ֆ���;Q)�B94�1�5�1-��`:�*kr_�Ō�<�Dke��]���5�B�V{����^���sm���?�J�"��:1�
�&����˷4���5��j"�eT2(S<]�]P�P)%bR\Yq��M��}��Zcw��|��o��/Ν;w2���PK7X/��ՕZ
g��իW�y�&W�^�,�z����~�ٴ��˒f1|���N1�`��Rĕ��FC������d�����b<U��G��J�JZOڞ��{�}ľ��w��}�D�D���g.����)�+ˍ?��`��YW~�Z�1�3,)ET��Z;�Є�[P��<.�`qe,�Cմ� ����~r��<�e��ke�Ln�YΔeiLW�e�I"�ꕽ�y|��L9�*
ߚ^4yU#�X�dR����EE��X���L&5o��ۿ�����Ν/i��c�
��v���T��\�����n�s��tL&���=�7��>�i
k�{h�%F%���Մ�܈��%�]�εk�p�Ѷ-�Ovx�����pn�g}	Ë�Az��㟷�J*I����������W���X��	�������%D�Y���[��3K�v���8A4�l.߿��x_�C π���U�a�x���}Z�3���{��&vټ�M����9 ��+\��a��j�M����� �㍎3��Y�)C���J�b$:�Ϟ�c�cK(˒<@�d2k�������9�?`4d����5�Ic�����[ܺu��W�������Gܹs��;Oh��Ҭe[c(�2�#�V��x�"��~�o_�(
�Y��M�Ǵ~�R!� A^A�9���j�3}ov8����=��nguss,����e�y�=�Nd?�U�K_%{�u���=���m����Z���.���4����z�ε�0Z�I�}ǹ�,�g>��8F���8W`l�ֈ�5�	��@��_�}�'���8��#$I�Ĩ��Q�ѨI��6a)vb��� u�>��B_i+ �S���&�<^��?=���m��wvA�J*¬��D�x������O̚@U��쀠`�a�q��[ܺ�[�(�I�<����|�)���S���`��QC�<X�X���Q)����*�X_�k�����/�՝<�W�]E�Y���t���a՟�ϼͫa��������S+��x8I3 s�`ur6s.u�������wr��<.��f���7�_s���v��'E�w�y��O!=+������7�#�d��ǴB_���cN2��O��%F�U���ZO�~������IX�-tL�v�M���Ο��Y��;�,�Wڑc=p�}��N<[��2>q'�I H�\?��7��z�K��)��x�^�[#��-6�礟S�T}V���f�g�2���Y�>�E�j��"�=�G�`>/�Zͯ����[f,!�ު�tm}��f��pΥ)����v�j��ε
ߢ����'PL���|���*�����}>|ȝ;w�]��SU�gQ+F��p=�L�ommq������u�666�L&|��W���?�w[!���tt� 1yF�7o���ߦ�*���r��]?~L]��f�\�����߆X�p�N���~�-H��y��=��޾�����ZyrtBx,�|F%���O��߅.^��~���=��n�>���Ua����[|�c��҆E�/��U����M��,�_g^�Ǖ��� �ˎ_�;�qΉsN�u��uZ�����������[_����O��G�7-F�VEE� ��r	�Y�}JJX^]�̩�+����}�n��'hBU��!e9�m2X[[���?�>|�ׯ_�ãG������/x��q���ɫ��Bm�^�o0�aL�h��͛7y��ﰹ��d2a{{��>������4�{�@U��6�"s�on���e���Y�d����X�L~�3kF{;������߱[��a�Dt��Iz��d����㣽��n҂e�N�!��g[�*�}��l���&A@���nU㉠�E�A���Y>Þ/�c�AO���~�o�?�	�y��q�Ӥb��eP'K��J�w��V����cL""�\a��1Xg���f�{.���;��g��ŵ<�%��Ր�GE����VTU5_i�1���
�f�F��v����8\�(�� ����&����G��7or��E��}>��s~��_�t{c�����$h�%З'����Wʲ��[����y��m6/l�t���`�����Oa��sߞ3}G��ۣ�^g9r���:�*�B��(_o������:H�Dn�t\ ��|�G�:"$zI�2"�������j&e��벤g��N���.tvϜ�%����2sܛY��+ow��'�Ó~}�ذ��>I>Б���2��S�����e_G,�w1;h�􄉱��9S:�ֈ�^ӌ���'�g?��Y���7(��������kn�E?�b"V���?���aޝ�B�Az��:?I�H�m�1�N�!�u�oB���o������;����ŋ�D?~ȧ�����/�~�F�*���ӗ�ж3���ck�"7n�`mm�m۲���xrH-�r�u��r츕ٷ-���8��g�o��W��93��m�Ukw,_kk^��<y�Ư׳��������g{����ѕ���u/<�f̋�N��%3��9�*��%��J���LO��=��;���<����q,�i�(���Eq��x����z��獛}���U+�Vމ�Κ5��5�����1gouߠ8[�ݢH	lJ�`,�d��|c)g�5�{�s8W�W�ٳσ�&3��^}���dp8��p.�ԂZ�p��%nݺŇ~ȕ+[���y��W_|ɝ/����!�� �ퟮs��|��������?��}�֥M���p�����rZ��x���m��M���c������� �\����X���z��"�x��BT>?h��$w�:��L�gX�W�<���3�)�F3S*Bf�̢�d���*�3�ǧ�O�J>(DMWh����J�m5�������~��p�5�Gu\���ī`�����^��ιcu½��/ɋN�2~��3}=��3} )%��.2�IuՕ�!�J_���/�E�g�g��
<�oz�	���|�.�n]c�4��5������@�����v,�8.���F�2/�7�t���\��1��Xm����p8dww��0�����f|����E~����e4z����~��U�i;cP�q��{\ڼ��H�6̚)��!�������]�dQ��%z֖ q\��i�h!�|��&n��8��K�z���>ޕ8���h�:�x��ǂ�[-�XT�0��^?�>��`�?~!(Q��,���*^���4��o�xn�����vL�1�9��@&溾�LW���@/<���7��5͋Ɏ�� p�ƋX��|?�}��3��2�{��nk��lB��Ĉ1QL(4�ʵ�����y��ę@�A�ɉU�D��"�d^�:)y�������u����z�*�������s�c]�]��bTK"֔T�u�p8��W��x�ob��`Pq��%޺z��]�^7��)�lK)�A��U��>�����_��_��w��`�x����';s��=�r���f?��f��:)��0b���q���Y��*qV& =�͸�N�xFW��
0����XT0ϋ����Ed�0'k��V6јȋ
5�=��~�Ȍkϼ��~��ǅ��9��90[a:�/�u;�wʉ�(����۷E�`0�,K'���Vq�)��y|�����q�����q��Ό�`�w7�ɈD1N[�$C`��r���{�3��ٺVZ��aJi�.���b4�{����2��_��'�bLs˓����yY�x��������ܾ}�����r��=�nr�)��*��[J4	Q!E!%�A�d˖6,,)$��|N�>W�Un�|(s5�&8����o�q�-�~���i3f����Y�|��OO�SwmI��~��
,L�v,*b�-r{&���������q����o�3��ߥ���TP�2�ޓ�Q̯�����:4�4E���}�]Q�l�_N8=/b5D�6ʲ�G)�:k��Y_��o[�FՀ�t�`�(
�4�(*Tc>>���!$R
�k��q����٬�mg��e*Wa
�GЀE���!N�X"�f�w�p8�mj��2�͘M'�豦�үB҅!oǀ�����%y��My��!׮]����?����u=/2��)%B�\K/g�?N�������|G�r�`+��:NwgN�W�uW��>�s���x߫�a�x�[. 9��{�Ngh�c�e�|!�е��DD�X+)E�օpoc��9%�-��i�fE�d���f)�&�Z�^D�r��Z���d�����۷y��	?����������"�7BϞ�Ч�\'@�H�!��	I��l�Rpue��?�ՔMl$�ّdH�`PJC���q��gO�9��#Ƙ���G��ٌ�F��⌥��X�4&�&R���!	�*�2�̍�B@K��A%a�+[QC�<p
T�+�d�`l�MCUX���/Ė���p��0&���P�:B:�.6_��A�#�,_(܀�j���W.1(]�ڰ����A�A�.P*)�"��#	V�,q�0k[|��x����d����F����t�C��p�2><d��C=~�ݯ�dg{�Է�R!�|��m|���{�_�N&=z4����<�GZ��k��}��܆�cY��鋗^^.k{����}�_�g
U�I�y���)�0)xx��b�ř@_;D��+*��;�a^b��%-m�.tƂu­���C�Ww�`{�EQ�������Kz�QG���&�������RV�M��W�^��$_Z�,n�UJߚRW������ɘ��`I+=<�������>m,�����6`lg���5�ѐ���J:�)�Õ�XT@c"��E�G�쀌���8ہD7}$�u1�� ���	!q��8�`I�����pPRV����䐃�]��'��|2�F�g�k��$��Z�ZT#I-��z�mnݾ��k7ؼ����pP�֕���iIE��4�.��*)F��Ě�l�C �@���T�ӥEQ ���T�m���Y=�+L�Ϧ�v�{�����d�`�z��2�t���O�}o_�������m�+,q?n�)��q�8
��_)��#����8fO櫲���{��y��V阽��E�ͳSG?��N1%IIŘ�ˈ��%�ŤP�&��s��-��߆�Od�׿;
�fC�j�>���8z#/?�t���{�q��E�������]����={�c��j5PUU�t���3�58�0z=N��L���oy�fm.�*������{�r]�4j�V��|ٳ~�q��I7hb0�@�E�ePٺ|�w�y�˗/�\���81����`'S8J�8�N��� &#*W`
Ga,�C��R�v�
+�Pƹ�bĊ �RXK+Î�2�W��1=ܣ�M��_�����3�ݽK�	c!)�W2鉭>������r��������K[����&
+�X'x���dM砪OU/�[[�����l>ى0�-X����Sȩ�r�ƈ��d��c���K&�CrEr���ު/�s㸔~ߝ'��q�ެ}����.zP�0��;��X�[8��yR�g��C�`(�b�Y�:����~	��Ԉ"��1u���Ι��<�aq&���j�J2h���Y���S�g���C�����6k������K���� �� �o�DoΜ+��Nu�    IDAT�~b�t��-ȀO��u�EG�gW뫃Mh b���ƐR�Z?C̳��E����:�~�cy5�� Y# �5�߼�����������¹��Y��0�m��ӿL�SЅ�����K;k�5�����93h�d=!BH�	p�r����e!(-)��+���3(+�z����������}m�C�؁"A�d0����[|������w�JH��{8��$c;p'���c{V=����wk��T!%Hm���&��,WR^�AE]�L��y�����$i�$�C�D9�����f����n�Xb�z x2pXf񀕖��鷾S�r���o~�����х²Fo����Ξ����>�{��)�Ŭ��󽐀F���ak��oz�q&��xo̚؂�u����E���X˫�eEJ���ڵklooc���*��)�锭�-��X�#�1��~�%!�Y0��������7e.� �~G!���I��D�8︐o�g�=]��9��2�e�Rg�c$a�8Z�;�}��?��ܼ�n7��-��&�0����w��$���~k���|Uf��ɶ�vђ@�#��2<7m5�� �QNhX ������dXMK�\�$�Q�U���s�#{������dVeuߪY�d�s�9'N���X�[���8KflB�C���`|~��?�c`D�T��1h��D��=](BU�)(	�u�%t*΂�w��!?��S�%�m�	�)�yۥګ��H�J�Đ�3�pr�>�l���ږu۰Y]��\a����)gGt];�],}uCUUx�ǂ��9�v�ۢ>�FXT3�K�,��ߴ�]~�fu���
���r�{��sr�.��,�Ec�Z?��9;A�D�u�İo�>j7E�4}��4# ���_�M��LGz���ϟ��y��@��T�=�g���@	U�mۑF0 ��V�?_��-h.3c7WWw����V����f٭z������3�EU�AS�2H�w���)��r��M��?���DY����/�3�2��j��A�&T���ВĚ�B?p�y�ܸD�0ҧ��$���B��Z��ڍ�����Ik,V�3]�wb4U6��ng��{c<<�*j���ܽ�wN��\A"���-�͆�=.�(�|��E�DM��.Z��'��ɳb�(xLヨg隖���eg�m�����ق��i�5!�d.2�g,Y�ʲ�,K�ީq81D��V�k�t<���6�e��X� i~Eeuu�'?�	?��_��ZQ��|�l��ݎ�n����iƍ�9��n���u��U��m�^������Ȭ��v�_^�ێ�m *�|ƃ{�y��#���������yA�X��HBL�(ߐ�t��~}�����4U6�߾����noo���2ӻS�~�y�c��(�1��nԑ�78���c�}�ѽŶ֎Ǹ�M��a-�1Fڪ�1�M|��wX��"�ҧm�g��ɒ����cdou��m�VUE�e4MCUU��.(˒�(���O�{�xæ�{���E��l0i;���'nR�7'�(�L��5�C&tB7��!!�q��Ǩʻ}ᛲkW��*�O�Ӭ��eYZP#�UΫ/y��%O�>e�^�c�\2����}H�գm{�lY����� �����v;b�cZ��:��I�SeWoi�5yn������?�Xi|U�!&�k���"�6�>R����(m�u���:ʲ�w��}��������3�2�*s\~��n7��*�2�����2qз��Ib��뢌,yq��8kH�����sN~�GGG\�ڂ��W��w> ���/��/~jbS�g�T�s(0�w����c���&�L	y�����l6c6���y�!�}�@fzb��X?$|� �Z�EQppp���"���%��_�6Қ�y����V�������l��e��l	a�FC�T25Q1� VL�$�F�l�/`��-�G�)��]��0��-�ŌˋWj2�db��M为��u�!�	��O�tp*�Hw}9�n���L�J�l�ح5�e�Պ�jQ	]�fĘ�֊�%=��a�!xBƔ��"D��;����m}�)&:����Q0�Md�k���#\�!MS�n9\츸�S������_��/{��"��Ξ�}�����ꞣ���@`l>0q��آm��)�G�T���l6�N
\~���.}tD��8>��3���M���"˩��3���9��T��Ѭb�
��c;f�3*>%^�	���Liw�t9���)���eH�t���D�03<�4#ֽ~�D�JG��iS��P���q��`�6��yEYΨ�/Y�~L\,���[�q��_=�i���-���R�O�D�Z��a$ �� _�ٚ�l��k�ը�ٗi޺%o΀|�N��e���Ƿ����so�o���ӣ#%`���"��c6��X,F	��븼��*��?ZyVrx�����NNNn|��޳�J����w��%����9�l���]N�RP�Y,c����^�FJ��������wI�<~��jQI[�.}ݬ"y��k�B�M��g����r)�ٷ�n��8o��jL��AEzd얛�@��G�T�s[�
��~������&�@��B��zE��HfY����nǫW�X.��y�l6c�^��hQ�F���cS�\G�M�pvvƿ�w?���ǜ���L�=�����{P%���C��I�)B47
5RAG��>��&3��:T��A#V�lh;���6^�z�j�����+�&vTT%�_C/^���v}���c�5j��	�?�,�ą��"��}e{��9���1�Rц���3d����?��l>�mClH�ж5�F��L�k.�/�;�[Q4M3r��|�]
-`�皻�K?�u�z������r9��<y2�?�٢k;88�v W+ EQpxxH�D�躖���1�$�4�ۮ�3G�ٔq(���2�q!Fc��1Ħ���:Z��ڭ�^��a���(��g�F�og �j��5F	�O�e9�U��O�Q����URu]ߨ��3l����T���1��u�͆�,_C ~{���m�
���c��gϞ��9�g/�!�����0�`��`"Q+�S����I�����91��V.z�`%K��%����h�c h���l�k:�`L�EQ7��5�5L:��b68}�MDd�V��7u����U����:ɹ��z$���d��63dY���1��y��[C^��yI���w��c7:|o�K}�����wk��g����T|xn�i����'�s�{�= qT_�z5�iV���@~ѿ�$u�!�%���,�'��!z�vsE�����bD�{�k3�&�6�=m���4eI�ACZo�Z�ױi�X҅���,{�Ӗ�Dxxg����wYU��tƒ��T���״&ݻwoD��-���!b���$�O�~�������n���n�b����HJ���M���iޯ��?�E��g�=�vOhۖ��3�;2�rK���x��W�&IC"���\z1�yyC[��܌�3�#��[�!���,�r��$�#�8g�rK���}�j�BO`z��a7���C~*=-f��,�XT)-�.!�m��5�> ���b�YƤkS�{����ϖ,���������3N_��nT�� Lc�o��eY�/{��%��1�Hc��4h��x��c:��N�8���j��}ey�>�I_�m��)]�m?�R�u�޽���GD1�gC�)5dYJ/�!��������� d����%��:x���	�W�{�5��j).
���������;��[o�r�N�68c��g���*1�[�H�~�P�sb�cg����־#���AlBp}M�ZK�&h}�\���V+b��e9:�������Y}gߜ����AJ��u�j��$��#f�� &B�l�:IKB��Dl/�# mDTq��ӴhD��p�<�)
�ҡ}1I�4|v�&�@�j|��f�Q�@mWՃ����yۊ���;������]�α\���}�sBӱ^�i뚮kGt�,Kf�YB�eH�����Pۓ�]�s���#�=zD�~��r~�v�����g-7Rh���;{�y�o
{LQc%���v���?��?#��f��
�<����ؓyz��ƨ���\B�CHE^�md��b���{�r�d>���l��j��wt�����	t���JK�F|װ�l��ի�^���jeڶ�U�1�"���ߴ�s��|�~�w7\]�����H�zo��ŝqR>>~��<~���7�?~<��?��c�裏n��<~������e�gv��a�QA�(j��w;ޑs.q�4N�p�T4L�餚���Ӷ�f<M�0\�N߳\.������|�ޚ��#Qގ�M�9Mͼs��y�"���b��w-�'�*��Q�ۤYB���GQ�HJ��Mڐy��?y~�PcZ�1��ƪ����rpp���)�|��NO	�ë%F����!t�\��؃[����::����\ڷa�{c��n����,���p��14�=��9UUqpp���!��h������5l�[�O��y���;w���rvv����&��%�J�e@�Ҽq߬S�M۔�2�wH�W�/�N��S�n�������l���Ÿ~ܤ8��=}(�@��8��n�_Z�25cb$�@�<p}?lgm�������W�5��2c9_pz�k3|�QgK���n|������y��v>�}�C�1���U]7��fS���Yu���V�������ݝ�鳏?���9|��G�������g������Ţ��=~�<~�8�'�m���u�e�������Ν;���ivQ��|����޽��������#��n��_�f�7���Ǯ[�_��?��r=�1�g���V�7��3�ϯ���.OO�Ν;������?��G������ӷ[�c�\z��0�p��(��Sq�����S��w���$N�3gpʦQ��Ѿ��n��e��'��T�,#�k=-#Bf�3�Y��2�K���]AL�!����	��Ȋg,wf��CUU l�k6�Mӌ�l6�ZKUU|�;����1��?�)?��QB�/m$�X��M\f!f�eNQdI�y�0i��.������9g�HS
9fdƎ�5�Z��1�W.c��sxx���]�,��
1���eM۶l6..V\^^��/�dl6>������y�=e1c�7c �x}f�Q�o�������`{�k���A�|>�9w#m;Eꦭ�Pձ�p<�1]ō�6#�eΠ}�zP'X����u�n�����ݎYYrtr¼�(r�s�*X.�{�=�+	��{���Xجa�3�����m�H�F��2�vm;8n��X�t�ģ��Є�;u�y��k��(�J��y/��$���h�����;��]8(�͂�My8߬����Y�i��E�m�����D���_�W�a��޺��f;��J8V;�{U����q	pڿn>��O���v'�[���Ƥ)�F����ٳ5����QY�f������w�Т�,�F �ЃI�]��֫PF]Gs$&�F#b�.�5�|�
�nr5}�J�h�0qI�,�vW����m��*)v;�c�U�pJ���C�u����#��>����sk��ιxvv�
�z�O:�R��h4�)�u�:��ؠw�����N^�IL��i�����������,˘�f8�n�o�F��}�q�\������kS�}P��T�������(����w��x��W�%˃��,�ˤ���|NUU��\�s~~�f�D�w�y��}�s��~�{��s>�O���3��Qr��V�^Ƈ4S�%���0:g_E��m68}��5���!��Jz�\Qi[�v[���Rf�jVb���9稪*��B��[�&İ$#xO�D�6�B�Gc���.��!�?�O��ǜ�]�HUUt݊B���f����&��w�E6� E1��5M3�]��ƈ���m[��-����|>MӼ6��E#���=X�4]�y�(�����G���{������#>|HY�����](�G�wPv��H�O�I4��Ū+=�_Ί��6Կ=��e�Uӡ�klB�ľ7�ZQ5ǉL�ƴ�Ĉq�U���(�5;1�V�.��F3+f'��,l4���D$X$8�A��UT�ݖ���HMl���hT5A4�5�v���fp�ҸZb�]yﵫ�0""b�����I�D]�z�g��%���:2o�ع�Bv���D�Js�p�!*�TH�M���K�F��f����fM�	Ar

�QP0N�yI�1I���9�s��U9���LͽJ�.S��Nb���Zڶ�9��J����=[����a������M��VN��ё�"��,DAMT�FUׇ݃ߵG��S?"y�KS$�3?�|��fLqu�'�_��5��?o�*+��kz��?��M��(�N�(o� d?�<=����FUӁo��E�ݝ�7���s~[��mc��ɞ�����3�#|	�-�kgJ(X_]1�9��9!��6\]mȲb��ʲ��|���]NNN��"��("4!�-(燨ɩ�m�qx�./_>��/���w����٫Wx�R��m��&�,�y�j�Z�?}�_1lR	Ŋ�3�!@����ޝy�Swqԥ�+����|�٤Pe�������]ץ���yY�u���"��(�˄��,G�py�e�kX�.���e�Г��o���Ֆ���@3Ќ��gcZm�b����.r$�<U�����%v���u�r?/g���̩��N�����N�������~�/׎H�n�%[��Z��x�#�y����� ��M��#%$�4���f@���������~����srr�Ç9::��@w:{y��t����Z�+�]�|���a��h�]�_^#���
11���FL��J��0b�11m���9uY�5Q�!Hf]$�Iʈ��� ���!�����3E�r�X���8��:&ؠѢ*�˽�]�dY^;��!�1b��ykmK:�`�M�mTTՅ]�cn6������	��jUc����D��ֹ����NUQQ�>�����i%5� jhDE�u��X[���:5]1�N���}�e;��Řh1�d�S���Ҫ��l��Ζ&���Wͮ�;;<�7�9�!�+3��u�e6k�j���������~�O�������5�o�@*Q��bT@}*ݠ@�I���.^ב���i����y�/B���T�'nH�"���Q�e��iï7u���OӖ"B��d8[�1�O#�%x� �A�\ˮlYg;|��
�g��W��@W̉\9Ǹ�g�Ny��W���6qآoA������1Ό±�9�.	['_������&��S�N�I��E$z��M�qxxȼ�06m�����n����kܮN�]V���'-Mo�\*r���W�����9����?����S�#��+���!�v����e�t*{P`��o�1Ӵ�4 ����o��:�y���c�n���!������ܽw��?>����|�ᇦm��ߋ/x��)/^�`�ZѶ-�k	a�:ٔ�*�$���ը��V�\�;s�Q�80*��x�J&J@�1�Vq QP��W�8���b��F���	^�rk�WBhQ��q	Ռ��n2K-֥�c�P�N�O��K���Y��5	~�C׷�T���}x}���m���Ö��*
EC$X�(�^�k0�͊�	A����2'�K���D4�BX7Ω�A�s�Q%FED""Qc4.˼F1�]�fm����La��f��k��<8yZh�c�w��3��umϲ,<���{�����������_��g"��r���rG�d�"�D���5Q}��N�0=�yD��?V}��u��7'ؾ�"���h�n*��6$e�#����۾Y���ĩ���O�����"_�l���X��"6-� �q��vӢq��6-�GK�,�f��>v��nP"B9�Q7���1����?pvz�v�P��w���� ��*(�GJ���ucRAI�:d�^$i����$ۍZZ�a���޽�F�e��f�P�%�K�'b�46k�@���X��Ҷ����s�뚑�:�?;�ɧ��{v|t��W�\^\�Q�?A����_���w����3��uh�o�L���4�3�7E�޴���!�5�J�4���;�-��?�GG�ѹL���cUU�m}V�Q��    IDATo��V+�?�ӧO9==e��"Q)\��D������Ԣ���Q;���+T��!*ɿC1Fz=M��Bc����з����j�9q�I�� ��	>`Ħn;�K뗵L�HU���1�nHE�&����±�w�J��1zBPp���*j�WY � E��@�j��XL�R�V��=�c��>!�"XcG�NH���HL���t����� �Gt����::�l�n��� b�GI7
C�X�GU$�2(�f�2���B���lV!F3�nU�s���ф��E�$�>{�������)����ݭ:r���uf�UjF�"����D��V�.���}K�µ0�t�o���C���������L�!��&���^�����42��T[K���,*P��E �@e��l������A#����@���#n1#���y�:�Ѿ3�Ř��9�S^�x���Wt��g�o8��̐;��\oi6M�v[|r�l����ٵ!�lL����}�o��9�s||�G?�pQQ�9���ټ�	�7+�%	}A�DM�I��ƞ�\Q�I��NB�EQ��S��� �H`����=��v[z�� �n�՛�~���?�toJ����Lm��,"c����>��C�����w��l��IloBTӶ����l����'=�a�z�S�����;���l"�b��R1�1���1!
1$�I�������1d�%�=�!ɤ%~VD�`\r$UQ�e�z�'��R�y�6��x]U%�y��\U�_�3Ϡ��0��u)#��<;�����۶��U�����`��%.'�]ZK��I��7�6�X,��QK�$�.l/�o��q�#���)H�#�Y�3 bDpVȲM�o��\���.#�G�;��NRp��Q�U���,���{Z�Z#�m���A�U��E�a��hu���+˟֮�������ӧ�[:}���j)")�TS�a��`H�nzw���+��_r��|����x����}�E��@D�O�����ЫwHߛ9��ocS����׶m����kG'�<z�}��>�Ō���2�ȋ
QC|�ֲ���5D�����8�XɈ�ӵ����W/h}ǃ{w��J���\UE�#�~_ץ��r��pq~I]��e�s��"�or�n8Q!@�c���~�*����C���!�������O?O)h���;��T9]w[ʲ�����y�3����w?`u���┋�s�֗d�cy0g�I���t��;{g_bӖk��=;Ӟ�S�ox̀N����5d���b>���������k��k�����t�3޷�Xʲd���牎�bS�D�P��mi�Ժ�w͘�v�Z4ڸyTET1�H�;�H�{G��A��W��(�'��[*����c�b��J:N�-�mI-!&D��_�D�5t����~t�Āok����it&�Q��?ט�®k'1F�bUN�<!v�TK�54J�:U�ś���8:"VA=�D�+0N� #DA%�XR����)�� X�I�u$��78k��tmHWbr��]K�Y֑4�u�6uhR�wl-bL:�oO��ɜ��Ǯ�|��I�y!�*bT����w�l�\)aU��s��r+�om�:@��,�����)G=���kT�!�����GNÄ3��k��-������<��S6���/�h�vTr��6]0~�׿������q�&Du���E�&�����8>L���ܻ�٬�{��1�.ru����n���1� ��$+`�`l���F�6Pf����.M�c^��+��^^D�4��l`躖�z�sx<EiF��� ��oZ�n��z����b�����<x���lF]�\\\pyy�u2rc$(h ��������'M��b�ɝ��*��O?��?������uMYe,����e�o䝳�m������q��=�{�f!���k��s��y2���s�ݻ�ݻw��Ί�ԫ�+��ù$�rqq������zX���Eǖ�0r�� �wF�	����9푿069� ����8�O��Ǻ����9@��e�	!v�~�!�{��:���@�u����@Q��5�O�FDL�H�9Bp=Zx���'�SJYBķ���x�1gm��r+1�H��!���&�`�D� ���1��D18��N!`A#���TH� "�9m����}.K��	tɡU�RA��)���c
:�4u��E���֊��k%7^M���/L���Q�u�uB�l[U���?��?2�J��_FUU,���TS����熿���q����.�}��#��Y$��$�v�t{��	��y�o����z��u�:1s���brH��~���y�	�w���T��\�k74�������@���=����X�E�`1�ٻι\����3�N_a�b�z�d�Źl,�0���dGׅ~&�/��u���c����}��Im	����n���+v�K|h0ɲ�5}Sy��Al��+˄V��Md����%WW�\\�%�2"w��a6/��¤#���;�~g�m�Uy�c6��Z��9���,�>}�ڸ��}�ћ~k�(�N���u�f��x�����L4�>C!�o78�]�h!/��~D�i4�E���2K)M��b{dӆ�'�T�Oȓ:))c!��	�A=��	�2V1�@��X0=�-e"ҹB��H܀��y�-�әQ=F!�*�IB �"!^#i`ȝE5��U�I�T$�J������Q^��Ū>C�������t�1H���}��ͮ{���5�K�֌���ǙaL��#y��|O�a_Je��з���H��ش��kE�����Jg��$D/Y���mp�ʖ!/Y�����:��<���5�}OU4�$���]#}İ����_w��& �O�������ސ�"���*��_��6ٴ
z��~]�0��ZF���@��lVr||ܣUk�f�fs�z����ݶy^bm�t�&E�=�Y�!:��i��*�(E&, v����ӗϙ�f=R��;c��'�f.Oܕ��ӵ1��L�;֙����q���+�>U�����������2�I��Jfe����w��O�h��̲Z�X.�TU�ԑe�횧Ϟpyy�'�|�j���'�����(R�|6+�w���:}?�9���X���~��Mg:�c�Z�l6��ݻ<z��}��k��ӷ>Ӡ�,˱��v�5+<x@��R������ *�H�ԗ� U%�^���`�s%#CA��%�D�����ñ�Z))%���(�Ӎ�؀s}#��WC���Dm����������'��W���i�����G�ff�Q ����%R�Qz~�D�I{p������{��m�
Ltt�?ǌ]� �$���\WYw��Y���E<��8��~��)�Z3:s��er�D`�X }�i�����?�8��EY�g�o�.���&��eծ(�:������ό��Y?�����ٟ�ٟ�.���J�ʕ�]�ԵA]Gɦ�r"��Ut1pqq��ppp����3��,�����7#�c����!�?��2�h�%�6�T�c:B�ݘ�S"���5�]�I�_�1=���M%ZTu�쫪��t� :�~��qkR���Q�9�W+�(����%.�8>>�Y5�C�����wPu�OgO�c�h�1Ĥ>ف.M~c0�al�n� �:�EL�䁮k�tI�uc:��̲↰��F��K�Ǜ��B=���BE1Z�S�i�bT8樷��`��eX�"��C���6,fs�Y���9�����k./ϰ�p�H���}�v[lY�-mӄ?<ZR��M����sv�WW���윧/�\�J��|A{��/W4u��Q�a;�qii�qBQt�c(ˊ]�b߀$O�����_{H�"��T�)�2U�)�Iʹ�'�4`5"�������5��N����]���ã9���E�'F!XG;���?��c|�l�5E�H᫳s��/ħ?��������n��a��k2�:�.8t;d�
�{�*�n:Z�Ĭ�n���G�*@�$D�د�W��:O3o�m���_.���Ͽ]�T�U��w��?����:Y;��h8;����o�#%��-&z�A�T2:brB�W[	X"&v=��}�,K���m��|��/^��,��ΑYG�8C�
�،�_����U��bA����1<z��|N�u���s������%���ylϰk����(�T�d�X���Z���+}���T��y�5[�U��!
��d����wԈo"�$U��H�q"i�	�����z7�A�92w���t��9�~����+f�*Q2d�&��@�Ћ��y��ډ)Ö�*� �'t�=��������_ЈnS�u�	�"�Nh��8�n�g�q��0M��7,Ĩ��WW����t7)*!]{Rv�ZK�K��&b5�������|kC��4�3b�X�����U�y��*ۧ�=��;���=�����r+���͑9�sng�e��7�?4ָ���bq������ܫr||�n��'?�	>('''��?��Ç|�;�[��ЦJ����f��>8'�A%r-r�����O�"���(�V+f����5a̶mS˜/5C��uUUq|rw��l��5�1de��b4�yvcQ��&UI6)�����4"�FޚI�J}z��K	��!��}&�]��6p=��sT���O�<��'ed�&n��Ʊ�D�e4�TM�׹a���cK2#��>����3^�xE�4x�l�B��������w�4���PM��Wu�SN����N��i����yV�>��qyy�RB:�$F�r>C$����~AA7�o;DW��PsN�v�<u�i�@��fGizD3"�6�a~��:���s���v|g�1%����D*�jO��:ƧGTԠ�;���Ħ=�m�)��(s��Q�A�y�ٰ�6��f��?E����}$i���ck�A��իWq��=���z̦
�r,�����M��6���qy�bWo��u�����9�>*1�^��5�RV�Y�o�njb���Y�(1�� kՈ�h�k��"j�ب�ֈ�tm�����.�� &b�11F%��Qɫ�'�1VĊ��%&�;l/�"Q�=�$�b�%&R,�ԀŰk�t�%�kɭ%K���m�c��#�!�M�PDERn]DDQcDȋ�!�:��V�h�ѐ�� ����$I���DMH�pbF���(z�F|[L����<ύB�#UQ�n6��ƽ:�l�3���Xt��^��f�uu�Ύ�Pxa�絬Vw�����>4��#w�]��Z,we�>]mοqy1__m���#r�.�͖O>���G~�_�:��[��~�������w����z�n�A�������c�!����u�{|ұy휦��s�7����c888������a���8�
�?R�;�IE>F�(�E���`$�/gE_u1.E$�7�dLS�)e.JP����װ6�C.+�6�kS
q$`kPZ���_��NSb7y	�>��zр�I2���'O>���Ã%��"��K<���#���c�ݎ���� J�yֻ���J"�����iȳ�!Jd�l�ϒ�rQlv�XU�/*��6�!�(��Sn�v���oB��3�����QV�jFQ$��#��A�+m͚t]c��a��u��imC�4dE��{��]��A^���Y{6��*q�G*�TO]�~�_�x�u��&�� �o�}�:1�����}u���LE{�A�����{1��!D%(X�1�r�9�����;	���ϟ��:!���z�}��^r#��0�^��NM�ӛ��m[��i��w�����GwX,c����fKV�D�]s�WWk�THB��qآ����A��^�Q5Zkk���ͮ �!Q�Zc%`�F#.�P�J�(i�S�F�� �ص�c0BT�h�E�ɜD��x�,��Q5	8%WL�Iu&����h��|L� �C�EoQE���C�ƣbS����'jp��bTo���Mu&����D5Q�(*&`Ԩ���^�DT����A%�:qV%D4L�����de~EP�ZŪQk�$�K^[P0Q��D�"����Z�}�pyV�l�n�?���ؼ��mk/W]4��ZSΗ/c>mB7��;5���ms�`S>}��r�f��ɬ)K[:g�u}L��ϖ������<���'���<����������~���<�麎��'�>�����z���:���uz��N�x����nJo��m�ޘ��}����X,������v��7:H{�Q�+�-�_�xfՒ�,8>>����fC�J拜��M��(g乣���,+0&�cL�Ve(�W�}$���e��-ƪ����[���q�y�˗�	[;�\��'H��p�wbBHZR���4u��O��η��-֤��(�4�6�����Ǯ�����$�@S�l�[ !�yVpxxؿޓg���<{���nGY���'�P䡿�~AE�1-L�˷�o߯!�r��}�/ƈW?��%)�Sf�;ܻw��|�^I{y�Q��a�|��{]��g4�ѣ1`p�����C�1�Vk�.׈���)���>�W��x���_�o�&"��篻��M��N���J����zA���j̐�����$g/�ɆÚ��ڶc)ˊ�G����|�;����=�����m9??�B��m^s��Nݾ�K����hc��Q�%�Yjƺ^�YoJ\Vp��{#��g�~���Ϲ�����紭��k|�gs�>�2#sE��U��,�X۱\΂�U\�bи���^Y�M����T7�1DDB�k'-5�0FZ�N{�R�bD��a��B�@�E�5�5�1#�%CU����Pi���AU� q�gD�H�C0�#ј$ *�l>����(��b�H!ΡN�LP�1�^@}J��֤�a4J��	"*B��Q�`� N�1"bzb���+`D,j��DL�1F��g8��N,N}aqI�P%KM݂�(Ɗ:�PE��'bTd���fWKS7��U��Qe���(��b��˳�6��6N�%&����]G��p���s�x������ӟ}2����Kg������~���{�71��gO������}�v�e�M�^�I����h�D�b5L~��Z�q��d������ hŵlF{�s粛|���A����������ײ�J����s��E��Lf��UE�%�n $j`�p0���x$�dO�T4�&6jJ���p�$��b���.����ͽ�t��`�}�7^4� �ɬ\���⶧�ͷ��ַn0M��@)�T->b��������.ZB�hm�T��+}�) A��(���ֈ�dD1ZU
4Zg,�e,��-m;�,�<xt��>��O�;Z�9��mFw~�2�G�a�m��Dƌ�(�x\���Ÿu�![Qr�y�eͣ����{�wSd1J�6��~���8����+{W�&��O�N��2V꬧!(|!����>x:��u��ǆ�A�0�%� xK�v�g̦�NC0jz!P"�$G*�	��{0���+��'�8<�zL�^ 2�E��2�H���4�?�'�'p�B�X,z��k�������Z��{~�q/<���v@��٘[�������+/�ҍk�l�@5�'�Gg.���m�6ı�8E"=?�u%��r���w�]i��<�gP�Q|����G�q����Ѡ�!u��>����k����1� ��D+��4@�_�&�"w&�m[;em3v��V���^�_B�6�(�\���>�Wo��V�g���Yk��+Wx�߿_ ܾ}[������Z��U�:(YԕX�ЎGE8���s�oo/���$(��tz �U5Q(
?j�6.di��ɲ�g��"`!4!�U"���ZP�NL�MJ��B�.Z' M�S*(+$�SBy��RBz/�tN� B�
1�/�`��2�XQ���B�P�F���gI0��R���)8�C0ʃBH!\�W�hB�Z��,=ai�.�M����BdƁ�o}pn[y�-�HJ���/��?F΅�y��;����_�B(u�>n��_�u��ڰ�f����2�����)^=?<���ի�x���������ʫׯ�����{�QU����5��M��Y,�H\�|�B�8�Z5U���J�I&� ��K���F�ןdu�P;-)D�o����J�_�.��9�~�u^}� �و�i��ڢ�sF����Ƶ����m��^"�    IDAT� *�B$8�d�s1��\ܬk��1�B�ՆJ�h]P/�@�#���ݽFg����c)�M�W��HV7"�
8p�&GQd���5��ªRQ5��%�t����X�4zW�Z+�Zi,	�zpF)�(��Ҷ�Q&��<�E{~&�1L�'N��1O�6@w���Ma���ה�EN%B�vL!X�*^�Qn��,�~�C}��(F�gG�h�����
�c��,/O'�����i�,�9���g)W��{��	����OJy������Y���_�����$?X�V�����X����]<FE�	R��d��ǝW�ɛ��;ܼv����іs�Y�q�ڵ�/n��|�����K�,˲��:ڄ��f\�������S/k���9|t�|�$7��tʍ�n�IE��`c�U��ٔ�h«�ޡm]�&����> Bt�t1>��/*����k�e+�:w���xY��g�TgR7�1b�_+���?�hƍ�r����]k�r~|,D��HQ��9���^-��΋�B�\V2m��cW�4���u�T"����)��-N1*8畲2H��W6x)�t��ޏ��FFI�*��J
�#��ҝ�,BK��I�U7¤V��A��R���U\�Q¨�DV�m��C��؂���5%����F{-D� ����+�Xu�C���<���uP�U��B@�&_��̜��if'�X��ű��+j�r��F�Vu�װƸ�mE���kN�3�PB0��6-c����@cãr��>��A�X,�G#����{�'2����2�̨�^��7�1�����?�?�z��M������X�i������,�������'Ҷm ̲��֯G9��'��l�N�?�#ȡد�'R1*��)�.�g�c4s����]��|>g<�!��F�1�;�ؖ���oq��mv�v{Ep�c�"���f��%8h��
�k-���UJe��q!2B"���{WnrkQ������}C��U���K��1[�X����ȁ�9�q�t�WcGJ	JS�%mk�.���A�<� (�̠���-��($BE��YI��
���Oi�$��e�/�VI�j��l^�x\��ƛ�� b͐�Q;�6���5�[�R��_i%vV�(YAH�X���ɶ!+[[[�y��������5��3�v<YW f�f�R�8E!E�۶e>��|ޯ-Ҝ�m��o�6�Vr�خSB��I���u�D��	�0���d��yԾl,m3����5����������F�&h�|���	����h�����b:����#|�}���)�{�"�3E1��O�� �m9:=c2��d@*���q1fk:cgo��x���uՀִHB�≕�A(���U�B��Y��A��Ω��_����:�3�te�e5,��$xӜ��4AklfDH)d�/��Zj���Ef����J���@��"ӍkE�&���a<��E��)R/3��v��j��Y�V���@.sh��Ω��ZZ�h\���-弆�	x��m0~�۶�ң��^kC�
�@�(*x�ڊ�P�IW*�t-���!����I�*���RZ��.SN���{�H���VZ�s�\ȫ��:hmCM.�R�;���0˰�b������ ȂZ[8�E봒N�����a��c�\:)�h�H��U���L_׳Ҷ���I���K��;�^{|�Xܽ{��J��G?�Q>�N3�n�\���rY���ٱ?��l�_�1j*W��_��)u����X.z~C�XQ�2M�E;;;��k^~�����<��h��4��HD��r	��y=O^��}�(Ek��ҥQ�aX#�h�h4ekk�K	[��QV�%�Ķ2EV d�m%M6�s,DId~;�]k,��Ź��ֱ-�{6u���"���qaPz���
�٬O5A_�f��ջ�HY��6�d:�!�+c:�,��ei0&��Ľ���n)�U��K��B�|�]4Yu��-&K�K�Sb	���*�?3�S��9pP�L�	����Ǉs#�>���n��,��0�8�r���n�x����Ŀ�d�w�L�� e���-n߾�1�b�c�X�����x�J� �{�(@/d)힎x���_Ş���W���"�08M�(놲�T����P�e���y�[,��|�f��b�7��f$=�yyv���H)���fgg�=�1>�ivv�z��ml��-�A�0�c<˘Lf��cw���-������z�eEU5̗͠i���ŕ���|o�ʃb�5���ն�vP�� ��(U���i�?��?�������cl�?��?6;wv�ݻ��ܽ{W�+�<�n������ �O���uM.��\	������t��6���ݻ]�6'�����׹�=���x�Aw�#���Wu��c����R�E&��t\�Z��w�����?.r9j��s����3ᔒ8ȥ�Rz�XN�B��.ŸiJi�N6۪�B�|ڢʕ��m_��p�p2/r�Î��K9�b\
�j4
EY�J� ��U= ��)�쁗R�u�hfM>�TB7e��,ggJim�k������'����ޘ�F����\iSN5��,F�O����������m;���G//���GcJ�+H�ܽ{W�����d0�a���r^~����'ׯ�����>0����-�,ʒ�|�U���M�s�jٮyI)
�@댋�9R(��":aܺ�{04䞥��1�:���0z5|]zm���E%���W1���Sc)�u��L%�Uu��/*&�	{{{��N�\�}/Ҷ-{y��,;���`�i���S��PJvi�mO;;�loo��k�`kg�E9G����ׯ_痿��ZK����o������X���mۧL��y��F�NJ�X�1������$:�$���R��D>����,K�g�ϳL�#B�8_��5e:����`��6F�mF��W=؊Q�؆-I!%�d=�������4ϴ����*Z����I��4Q�l8��s��z�F1.2Dp|���<|������_�¨JȾ��t�s�\L��0�IU-���f:�0�a>?gR�}1E����%���B�P&R���ӚϺ~�⡽��l����阓cz�t�P�uEX�������G9]������ �4���.:��PUι^�nx^J���";U��c�ұ��k0�B)�K����4���E�W%R����svr�������7پ��:fY�F�ؼ��>����`r4�a�����O�1,�U_����˪{�h\�ل��bL�:>��I�����ߋ� BD�����j:۲U]����Z�N-����]�����O�n�S�4h{�O��O�B�w���@�v/ ��Y�ON3�d��u����������~��B�&=��m��+���������w�>����+ ~�_��O�I,����],�)�O~�Ez�}��������L:�&*��O��Z�{>�������&��𘦶\,TU��m�;⻖Q�$6�o��|�����kO�mگ�n����Sۜ��	C��&l�� V��H�nBNN����ϱ6�����9:�(��l���6�ٌ�h��2�R,�K�m�P�5��ؑAJ�Σ��ry�w-R�.*�N"�lo]�ڵk(ex3�,�"���׫v������o$��1%�V��R��r�����Bj�#:N��zK]5ض霅�P;nd�g�e<)�(���K׹ru�,����d���y�8���
NRt,�x��k��;<ݵ�a��%i�]8R����cGGG�����7��|��(-E?߅ E�dq.���>(|�B���_�E>��
]�Pֹ��]�>ϲ�R����v��5�N��Y����&��4PI�V���Ǯ
�E�s��+_�KW@V)��CXkeY�<���ixmdX�nױ��#�Jc1���,��w6��9#��"���T�1|>}��a�.!��j���%:�v����\\,8?��kAz]��Z�������y�|hl0:ڹ ���8/���_�n�W�~@�W�$!�B����֜R���-F���%�V���1.+���B5ֲ\V]��AL�@�GLR4 .�q�{��;�Х�:5!e�_�S ��FA��{��D�u2�����_l��%1�+�)���,�Ƈ�׋q���R6Q|��M��Fi��He]!����a���=�HK�u�tE�E�G)cd*h���J��/�~��n���x�=ί���s�]��@��$>�F	���qH�2����<x�����s� :��ὥi,�q�2B!�Qp��0N��0��(2ʺ�:��b�G/,� ��qL�&�(��]�$��b�/����>��s`�s!m:m�2?�`~~A]V�F�ј�Hk�u՝k�c�Z�4-��<Q�5˺BJ:0+x�]����Ż�������_w��߄םM������5m��@��C��/�����#|��E)Z���!��Tb6F�2��z:~���] 9 p��o�RA�R��i�
! ���T��s4�C�6ri۶����~s�F��OT����'���:3��BPwm���$�_�٬�gi[��%U�62��U:����J��"�`�Rʠ��� ��r#+����}/g/�͸�A�*쎔z�;ޮ.�j�[��L+#�m+�Hmc����������lş��DN�[�l����I�䋤��퐿�*��b��~���փ�T��-;u]����5��x��A�Q�͒�ىo��ki����L_���x!�"D�hO��-	�&��E����c��l_٢�� VU�_�H<�L���bY ��u�x}%��9QH�-����Z"�Ƈ��A'�#�z�T���-R	��<2�6EⳮsN���{R��E->(�Δn��v��0ґ����&�֚<���۷oRU�pzzJ�ƴ���IN�2nܸ�h4�������DG��� ���N�`�S�C:F����Ն@-X�C���k���4��}l}:�����f�Kkݧ8S����UJQ5yV :�<:F���YA��H�P]z�B�tp��^?��2��>��-���N�B�H-�
�����n.|X�9���t,�
�aT3=��J�h��&�7=��)%]���|�|�<�i�lL\o�~J�a#0M=uE,8�b����� �B�B �]�7��_�	��F�Aߏ~����VB���k�Dx�\��M��=��r_�QMc�VBi���	��������,k�]!GU�4sXq�I�O���G�@�u���@_��z�=/�K��fD#mr)�eQ~"�z�`a�֚z (�x۠��f~qF]��#9wTh�rk�t���"dL��`l�-K�����N��Y����ՂE9�n+���X-�k8���_F�R�\�0W�ù(vj�AI�:���}l�����،<�jg��w9*ʾ��Z�����=v�jI���`��ԇX�m��M;���"I�Em �}#���j���#¡K��o ������tʝ[���%�lo��3�Q#D�f��7n�e�>���������n��R�i^��|���xM�9̗��Cp�����ۜ�B�\nC��#
<��k�ް7y_������ZO�bb�4�d�QD�*��*���يk����f�A/���E��#GXE�D !Bt���*��!F�Et&����ԋ<��t�����Ɇ�z��4�ctUB,KiݢXU�6�W�~Ew��ή�����>:G���7"/�pa�r��Ʌ_�WԞ����?V��Z�L�Z_�PI�}�loX/F���!h��Bʖ�jp6V<�e�b�`�\R՝j�`���gll��GEV�6A��ؐ��;������nO�����i#}����HBFmom��=��~d�8P�Kc����bR�T� c�B�ض�#��n,ZOb@Į�6�M`Q-�M��W�%ی��Q���۟됬�eYWuk�wR+��նu(�P�'ޢ�D�碦_��v�z�.��c�g�/5tH6������ �����(� 6\�s���d?�g����lm��ٙ"$�&S�� XJ�u[��LF�Q��� o-Ai:l�G�DQ��:ܠsI�δQ��˾�%�>R�v��xX���@k�^d��=+z��J`��[�	!8??,0��%�p;	��<��{�W^����N�^k&�(g"%k�����A���`�\������w���i�}���k���/t�͡�v��m*lS�J��º��u�2'{�;j��s3���M��a�_j����>��|�9�v�AV?��c��N1B���]1�s�{'D����E&�pA��?Uw��w����ϔ���i���K/�d\��ڦ�i�ۡ�oi����1�MdB(B`�����CU�,�Kʲ�i�ޫ��L<y<��|��RR$.ti�4!C���K��~ÈFz���5ӂ7��t7��K3D�	�u�5Z!B����M�S��6ѳ�]�^A���m� d�<�9��6t���bU�`p�%�g(=[Z���]����^>�^k����09L������%�R ��?�w��9�[���g��l�z���k+����Jhvw�0�ls~�����z�!���b��m�@a�jx�C`ӟS�u�����'�c�|So�����
@�llϩ���{7�1���w��Z�CL��h����G�M���	e��;��u�����Zں�>?g2ʘ��\\��qqq�����8��iKU̻��ܹs��7o2�N{�����J�����G�qxx�GĆ��i6��Y�q��-^�u���h۶�qxx�9L�OgyT�t!T�'&�-��*�����ʕ+loψ}������dru�9��!��߿߯ǩ:XJ�Gע|�YbZ4�@�,MS�45F\���՘N���4�W�<U�.պN�H�~e�������}�C)���	K��&�)rYe�g7�v��<���  ����',�K)�T!��)������e���!{&����Ea��B�.��M����ŭ��!d.�Y�ڶM�P5�Wl�4\\\pvv�"��{z<���a�b�e�͎+/h)�>L�$]�M�aU`\��?p��TBpx�ҴqS2]�!.Tݿ������RH���xD�F����Wd��Z���ֶ����9εa�F��Ǐ���REj:ס7/���d����{\��G9��]�"���=����X�� ���Ǳ�(&�|�\�r�G���s||�Ėa�'�6��#+_�ml�������z����*��}��� EH2u�I��X�y��}�1����y5M#[ư\�,�
�$����(u^r�:����=><�(88�k�"�D���d���-i����|�����7�d{{���^$�/�ܿ�w�}�>����}���Z���lM�N������?����e���>�������=g3����&r�V�h�x<�ڵkloﲻ{��l�U[�uG*��6!B�Fݤ��L�yN�\a�!�/Yn4-�֦}�Ź����=�6#�J���x=7��%o���=���E�}��5]���22����{��%�u��g�Dk[��D�TȂ�)�wNxB�k�����X��'?�r{H_ۯ͞�*���ۚ��Bη��(������C�~{g�:[�mB�z�y�E����t���#����JM��Y�e����u֥Z��fк���NF�U�}3B2�`]����)�#P*0�Bȼ����2��N@+R{-O� H�!r�\@���Œ�j�"�;�"�׫���=��#�ж+1X����N��B#��X�AZpb��;hs��\ń	�Y�-1£q=A^"A��;!��b��"����Ł�ӿ��T�W@ ױSIE�5����,>�m^�l^st���6�RKPc��tdN2��A��l���.g瞳������;�!M�rxx�T�(�4
)A����Z�l�2�Rh$���8�dΣZK)v���b
�G��GT�#\3c>o�׊2LX�#=N7�� L�h�/tu���ʣĂ�{���������	/����#>�茪�bUMۖ]1��i���S�F���A�!	,|p�#>��N��ͮI�1ʵ0Q�i�αl�����Z�Lf����    IDAT�r=XQ�l�����a[a/.x��}�|��5|��G=�mK\��"$�o�^�oα����(�>�����!o����(]����t�W9e�
��h��#�2
�y�o3����_��w�-����_B�d�s�&к@���AP7'y6��+���0�����{�G���y��QL����¤�c����O��ã{d��)Y��i�[��	�;Zo1�m|0\�im9)+�|IiA�]\�chj�4[ܣ�-�y�#���-M�E�����O??���9���x K���K�+32���~YU���HtW���Q���Zl� dF��ف�ʠZZ	��u�[]�%��p_J�Q�d2YE���W��L�3�`�$؊Q����Z���m��]�gu�PE+����'~���5��v���O~�g���F���e�������m4��mS�m���qV�\ۚ�r1�"!hk�H�ZY������t��S}2��i���<~��'m:�M��I\�gِ?L$sί���+%k �@7��--"��I��e�����ަ���8Kq\���pzz���9��"�r�_�o�w�R�[[[L&ڶ���,VC�RA�-u]�eLM��]pzz
�����t� �F�u9�1)
����0jZ���c�2X�%��R�bDEM[u�4��9??���ggg�(t@
�)�e>,UU�ӟ����^��������^A$���\�� �Eɣ�c�j%>�9�6��Y��_�6]���1J����*I)�N�YN]�#���>���G9���|�"�D�n[�f������(i�9�~x�G�c�Y$��UJ!t�����9;;�W_����=�����ƭ[�\����"�
�����ߡiJ��k���=���lW*�aEt����޵\�ٍ�����&�=�;WؙL�'/���n8<<���}���p���b�������et��O�~}�1��dC�4����&��2��g�&�h���v~}�4������<?�=��lD�N!��cc@�	)����Tq�w�{�m[?Q�|��ھR�D��o��y�P���������>����y�|欕)%�8��2��I�uC�Y�n��?ib=m�]69�mN���0��<�g|��6�7\��0!�m�I�V����1i��X�f�{��sH��z�*����P'��x�ˈ$!�?����}�������I�t�fdQ�,�cggg�����>GG'�Ŝb�Q6U�Df��޺��JF��8M�s0�C+�4�}C�<��P�������9:9������R��ô/ҵ�ƴ�!����Q/K�}��-B���� ��K�p�tk2��o}�;�nvU����s��d{{�k׮E���'g�<x���t!�����4K �����~CmMc�n�m�_ҡ,�`6�f<���t8�y�`������cL�۶�J1.F\ݺ��{�Ř��өb�&�)gg�|Y#��
.��he@)������|�{�����s��U�Q1c
�� I11�~U#��(m����()P�T� ��,�|��'����f3�2(�3ݽwx�o�Z��Ԓ�(�m�g�~�/~��}�q}.ж5�iim���E	I��]˦S�i��� ��5�`����mF�6�线4X9KB���)�����Cǉ}���?�������f1x!;�2!@�y��|�h۶m�.���eO���y�PJ��u���������U�^�u%�i���n�z���3�c�/��I���?)�&�����z�M�˵�ަ'�����=�t�B�����$�O�(wQu'j��V��<�#}�i�=�}�-��C���^�@���0��w����"�z�m�`%��$�?����i��T�����:23��.��f�j���"��j�Nx���6�4��9�E.��0�B�0�I-τ�Zj�.]�,U=_E<dlٖ��>D����j��E9?���u���3<x�Ғ�r���)�����C�b��7�z�:��'a�)�Z+��7\��4�֪`���,�x��Ke�{�TdZ�n������W��/x��88���&G�8}kɌbR����~HӾʕ+c�f��x�W��u��ѽO8�#@�LNn��X/OGl�v���m^z�6W�^�+�r���m\g�D
M�%���w�޴-6x~��_�����xo�ʐ	�ف�����T�9!������l^���j�NNN��_�����?e����;/R,�����p�F�n�t��)�r�7#zC����a�m���y���ק��/�qY�am����sx���ވ.
!�A�����|�*���w��]N�|m_�.}?��G�,)G�r��<7�}k�"ǅ<X[�U�ؾ��m���n5���+B?	����`6'³#}���gġm
i�k�T���&hn�����3-v�h�"�i��7�҂��qn7���'�����)�KH�ٞL���6̛�
��TfB�{���I�%�E��/��<�p��������)Zo���KKY��pq���I<�'�g�<Rx$�Jx�z�s-UY"���Ѻ�T���G����nh��E=%#J�����cQ�?:��.b��!k���2s�_֑̿����������Q*� ]��1�!p��M�wv����{N��D]6�i�g��xo���Z�@��-e���K-�����Dmȶn�R�<��9?��ˇ�>�v���@l��#׆"74����|�U��aRL1f��Uv��"��X+^�4��A*�����[������Ɉl�̜����G�89����n��׸ze�"����o��Q���S>�A�Hap>�Enȵ��Nb�*99:`<���������-���}�O�	�Qt�5�9��E=���#x�Qp�Y%����˂CG/9C'p3�;�5x�|��eA�V�Li�Rq�w\�ZO�򑻙���� �y�k2!��!��}�i/..��/���E��I�>U���fu!��.>��=��R8�2k]�"y�A�tΒw�Ti,�G�6A�����'�U/� ���'�Uz���n�06m<��u6\L�����M��t��ӳi�s��9���@��@����0��#i�)J�e#cG�t�����soC�{��(��>V޸q�o������IPU�Vv������#���� �7�.(��3��F
��l@k�eTu��);�>�(f��k�LJ2[
��)�@����)���T��ց�vR���˷��-B���lmm1G�7�N�������D�.wP�|2f�6l��MkЗݒ�L]V�4�b�����hIP� =���P�������2����Lg�Qڠ�F�����G\�q�7��m�����;c���9����+�������!3���)o~�[ 3�v�dň�_�;�1ϸ��<��n�Jl"���r*DY�kj+�]KSW�u	�#e�ZVZ�L�ZK�mc�8HB����ȠR���:��63J	lmfAV�T�&ْ��Pӵi�����w��a���;��瓢|�<BH����(*� ���]q` ��T��/���9B_�W�}o��vѶ���#��*����Rd��s�;'���d˪�5��R Ն��:�2�7�'EF�'z��ϻ�Ƕy<���_Ԟ�"H^�Uc��_������{~<GÁ7�?6��.Z����>k[��b�m�l'�b[��}J$�U7����k�x2����h���Oxh[�/N��BjW��˯F}�N,7����CzK[/pv̸�L'�MC�ZH�-}A��(+ٽ}qԧd�

.~^��l_A/�,D'D��\�޴iꔢ+�G��ҭ[\�~�����6lmm��=������C>��s>��3���d��R�9PisY�����:g�!1�&�b�O?/|_к�-�Z��#��<S4�pX�"���.�������}˻��:Y�ڠ��z�:CX����;�����?�6W�_�0����'���|��y����G|��4U���n��c<�p���L�S��#ڟ����#��drL$�E���6Ff�%3D'��%���K�H|yD�*�S�&�s�ZE����/��G�9��^�o0��Q�˲O_��n�����@��>����JC:A��د7�!RI%ʵNz��!���l�/tB_�W�}Y�����N��`~h��V��Xj�#B|P���\\�b������ڶ�ҽr����j��\О����_�'�Ӣ|O����MI�.W `��6mC�Q1�.=��=�mr�.��<��y�n�U%o�e���]B`�D��޵έ]��jrP�g�EH0&c:����KU׼���\0�M�_q��+\�v���=��������R�������'L��'��e�s��N�?BG1��zįA�nu\2F���ƬG�AU!�`�V��D�SO��0�DG��U�����:�m�N�r||�2v����ˊ�j(�&�d�b>_P�j��������zd��q����i�T��� |C���%A*>�
���e	�cr���	�~~���9�o]#�69٨��k�|L�O�fʝW��|����=����:��䀏?|�w��w��3*&h3bY9��'ܫlӐ��ֈQ1�(
2}��ͽ�?���1AI��8��5��:���#eҿ��a��a{�T��[,bˌ�}�m)�k׶4my���;�w��	\]f鵛���Vlϲ��!)36�	�9�.=�'�כ�/t��Y�"���
�۶�vޣ��(��J[�6~���EQ!�L��[���·+�h!����9+ j=���Ӯ����p�X�QC	V��4d����~�EC`�xp J�~�%��m��S
�o�tC�LmZz,�K�RvZ������g%��������A|�^j�7Y#D�3��z~IU-㢗�]�2��\�w��	��A�:��$���J�`mۢ�^S�-��@�����W=#��燭�ڶ[ػ��m�RQ��...PJQ��r�7t�x.�%�~�m	��V��ӽI"�1��y�.p�����Y���"j��lw�t�ŽO>�O>A�N�΅���P=??G�t:f�5鮅Z��q�	��xa"N��x��8,�HU�����Ti�e87攎�R3M��ܼy�s��atN���%�~�9�Ucx��7�&����,%�ɬ�F�e�d4��D�X��|K�$�eS�yF��(�춉�i��j�B0Oh��O�E�G�G�@�#�K���$�P�5����!(�b��3&�)��S׎�7n�ƛ�ag�!X�Q�x�d��?x��G��#S#�o�1�L�8?��'q��o�v�I�G 0o*�]��믿�{}���D�ڶ��]d`-!8��h�=�}w���"G"��e�
i����MS�ܬҠ1z[\>+/i���Ul��/��D�e����f�Wi]��Eֆ�9Yz<��9}�����&�iHQH�6�M)�Z��dY���jq���G!��#2���Z�P���t~t�:�����dk�oZ�Fk-�.r���͵{�ry� ʇ@�C|6+�`5���L�o剈u�1�w����O�e��
�o�f�ox�c�*웑���!��;'�I�����t���]��\��7a�]�a�Lj����5Z�l=��&�����w5nW�b� �Ĳc����)3��lo���͛�<ċ�h�sx���~�s�O�;����3�A�B�9 ���)걊\���}!���9o�c�2�qcy���|�7n��g��͛�w���	�n޼ɭ[/���e�zf��8L�{�c�E�%s��n1Ҵrpc$�XI- \��'b�G�G��cB
�A�h�L��B�T��#
d"V�m�x��u�'̗%J��b���t̍�7�y���%! e�ֵ?!�'bJ�!E�:e�+� +P4�Ц5<i�^���q6�6���(CN�e���|2��S��c��K��9��|:.�c$4�5�S}p��,)�����5���F�CX�Z�f&��[o�~�<������������n<��&�����Jd�û�!a�����ZOUU}��չ��5�N�%���$�#V�ڢ�eY/߰\./%s@�	�6%W��>zR�q�zuB���wi߫W���&ppp�sm����s�{�1�F�~[�oӫ^'���6E)ʴj����m܊���;�N��൑��X�9Ej�dy���yUrpp@Ӷ��#~�o�u,l0
k�Rj�2��������+��L&���7�:����<v�H}WS�7i"<{ %෪��w�v/�T�l�M���C...��f\�~���6U���_���l6coo����_�����-�n_����'8��m���XW�����.8l��@J���:"j�I�q��k �Z#�J�,� �֝p�H�Q2�輏�`	�fgg��~�����1_�� i��m$�h��h�k׮��K�����-��(�8օҤH1D �틄�,�c  �߀��W�MD���k_�Ս��_��۳��X~���\]�gR6�POs�7���a��y�e��!(�cr
c���Z��8F��b�M�I!*˼Tm^
{��6��N�Aߵk�dQUҵm!
�mx	P�����&?�%W���ٝ�{>FD�SD&3IV�J]��%Ah@���� �hh)�J�6h!h���$�����Ph4��"����$YIfdL>��fv��{���##��,�ٴ����xG��|�;�q V�ng!�Ty:���V�N�q��"lӃW7f��.rڽ��`a�:)���ӿE�J�Q��?W�����
�?L*C��:\-����͛7{q�rqqA]����_���~���?�n�d|�M�}
���c�o=S7�j���-���s
�v'�!��u�,�8::��F���E�ц���s�3���py��~�9M�k�&�US�i������_��_SE^Q�K��of,����k ���/q*~0��������y��	�����w�]�x�.W��]Ĺ���d�ܦ4UU�u}��1-�َ����c��U��� @�F�"%�^���_�d>M�l��1Ɓz���FR@5����X�'-x�iRpt|���w��Z�� � %vr�|FQ8#����Vc7�`�Ez��S���i=�Ȁ�+=�A�b�%����1FT�L�!����^sJ@<��!�X�D�jp>���N?g��+�p�Z6|��w?wwN���S�]��]���e�����bY�V�1"��k!�x�
���8F���Gu���_��?*l��������hT��2�!�6u��M3�<��@�Ո=���y㺛lhV=M+�P�e�NlW��:-�ˀ��Ŵ@�Ĥ��tLA�"��f���i�X��B_��w۟籧��1�ئ�v [y��Z���)��P�+�v��x!�~�>7};�=���+l���4-��~��|�;X���ϸl\f(\IY��tng�o��&�~�9��4MC���0����t����4�����U����.1�7`��϶��}�����l�S9�T���Y��uC���s~�ӟ1+g�G��b�prr£G���@2f��WdW�]�}zs*ȏ=K6ݗ�N��-�q��&*��v+���5�w�}�b�%���fB*�Qk32���ɞ�e��4g��rA] $�؂���Ѕҹ��_�X�f�%�!�%�;��3 *1.Ukƹ�uC��|����8�y/��@��n ��j���_���]��)�����Q`���l6)/�q[@�2�AMU��i,��u�@|�_{#?~'���=�������;+�2^\�1bct!҃�8.�S[��؀i��*����ލ�v���D�RNۮ C��f��`L?{��/�������_��]a� (�����o�Y,���^�S5d�
��θ.��c��
���������<Ϲ�����t|�(�Y��X@x'��ٕ>�4���3��!}2�]�e��ߧ���}��o����_���ڶe�ڑqN�m
��4?��OY,<=9�k#m�	!�����;�|�q�M���/*�~`ڧL���~:ޏ��r��g    IDAT���x��	�}����T����_>�����9�����o�W�B�qxlH��뒗�`uc�h���'
�k\@�C	
��z���s�L2ж>z�lBǦ��1DI�W1�z�e0)�,��jr6lښB3�v�A�jE���_Ij?*x]NZ���a;g��w�Ok?����1����Ϝ��o��F4��]�igN��]V�y�^���]���_zc�G"PU{�<������Vk��?��˲*���
	�*�JQ	Ƙ׸n��������,�[�.����m+H$�Du�*���T�0�`�Y@w�5��l\���2r�:�D�����rd�՝�q��M�_|���a�ڶM��5�H���m0Nd�
Y�.h�0j_�~�/�x���]�ї���������_'��y���i��, �l^H�W^6~�v�@������[�U��{�ɓ'H/#���O��|����٬��2���&����#BE��%������O?;�Ó�G���/.iZ߳'��נI�f�+�(ڂ����\0�&'��j���10��|�Ij���P�%1��"'ONyzr�r���|NPX�j��dY*�I��  s��$ ����!JL���d�w�o�AVfUNV䈳h��+}��՟!���OQ��,[�B�e�QSg��1�N���^9?_�\%V��cFr��i��3�.3�J��,Q�.D2 uߵ��M@�v-�}fZ@,�f�,I�����B ���#2^������Cfh7�m?�i��1ﶰ���u߱�ױ�S"c�=�}q�����o�믿����׿�m�"BQ��Z�AИGW��ߏ�j��裏����Z��bv�W�q���B����a��M|�Dc u�<v�������U�o�u���N-[�y����:�su[_��&�aBiۖ���T�>{��������l�����|���ݞ���}�睛��Ƙd��4�8���W�s؍��k���|>�/�O�>e6��;w��?�c*�|��gt�S�9���*�M������/	�_ �Յ�m[...x�p���%u�����5�>�]�]������:��-QO[��.`]�Q��(�h�~��d������A��k3ʪ��o���]@>0.۟�4���k�P�=HR�e
�F�����d����([����&�Xr�&�&���_���<x���kpE�s9�1-U^2�U�U���1�_;bo/��9�+0���gR������Y��X��m[�������h�2}�=����̐)��i����o����>,^����#9U�c�Z��\�8<���o����w����m�K�~���\o�!�<�؈1?}�C���;8�����r���zï����j_W���<c�*�͆.���p�f��&���!G�`����7H�%K�A׶�8�������G�tL7XY�}9}���%ٗ8���� ��{x]Zvxn�����kw+la��4(��g��:i�h:Ď;�����1��Q��#6st"C�E��!�}�%���������L�b�f[��������%fk��4eq԰�g��ĎE��9��=!�(��?�I{�؝�v�� ����m[�>}:�F�g�`�1�F�:1�"�` ���H9[`l�f��X3�-�B��d�h�1l0����,^-j0J�5��ir��oY>=�,�4���~����}�EG�C����f�SBlh|�j�A�/����J&�e�/@
px�k��ڂ<? R�v�ɖ/u��7�^b\A�AME�w����,Ѯ�v-�2��A������f��g���~9ccN��9�+�l�D����%ưI��,�ܤ�0�1�brCk4Z�1ڦ���nr����bFפ GE��s�_���:�񂱞M��5�r���KU?@��<_|�>o�(6�>�l@�
��p��&Ȝ�7XSp�v�0�Ő�!(��D����φr�2+�v	�ѵ3j_�X��7��	��%F#y�g�>������'?ͪn�\�
(Lj�+�d�x�6o�s��|�����#��32W��!M$�>uGQO�"��
��hP��2a�˜�)MS��[�IZ���s8OC�Q�C�?C�>O�r�}%�
�:�d�b���IZ���d��to�|��>���|�,�z��<�ɭ#DM�(>��A�1�4M�E}��za�WEE��mOz}�z�K�fgq6I��2���uڶ�j����߼���|�?�����>{�����&s�����ͦ�+3��6t"񍯾z?~W�8la/�ce�|�FD�#�aA"���X�׉i�!�Eۚ��x핅R�EU�,3��JQ���Ij���O���اo����=�}�ݸñxј��#�m��دM#�ADݶ�4����G������u����E�/ұL����x�v�M ܾ6U�]}�0���W\_	=��k��9����Y�H}?SjS�퀚�ӅK��=� 2���y*�@���^�7��5j_��} 40��u��Q��,P���oB���P1� E�%��j�P٫22"��s|S��Yb�B�A'��5=���[Ӹ�=S5���c! A12�=���� b88ا����4vm��eܸ�*��������=��v�%ӂ��|�D�F%�U�K�K�["�.Y�Q��])Y8Ǭ,	]�z��,*Y��S�k�CQ� X�vM�58gp���}J ����M[?����b��n��;�?�=��&Fx������֍~��ۥ��eb�h�I��]��ד6\7�O������A�\S���\2 �ymZ�7�[_5�:����[���g5b1��ɡ9���Q�����7o�^{�����tE��˽�m�\_,�e6_/�U3�F��S#�]��߷}��oZ�����<�YQ�m��ں ����""��L�5��z��TkS�5�B�P�Fa6�spp���UUa����d��7��h�	;U��1[�U��&�]��U���tz��ƴ���s�D �l���=�Z�(��dw{���դI|��@z`���Ƌ�PI�{췟5�tL�8��ɳ�Ƨ��Ŝyf!�t�s�ӄ��D��	��:���*1�����CKQmϑ�#���Lc� &��o��Mz%VU�7c�����7߸����g�Y-ϒ�N,m���\�+'/��DC�$��{8�����oq��c��%��s�^�xM���.Ϙ-�S��$��yU�g�^�k�T���&}ڬ�ǿ��0�z}�����,�)���r���������#n�~��܁n�я��:��A�a�����7��Fb��	��J& ���4�b��%�EA����A4���;�dF��5��5upq�����`��uZ��"���Dv��a]�������$���+�͒��CL0Wҟ��cj��1q	p:�(�kDl���+��WOJ_o>�.��ʀ��D�����(} p��iX�ZxMר�m���AS;df�4n�2�޳W�Q�mӐK�yꮥ(
n�r��w���l��?��}���;˪�m��z��iV����xs1�F,D�R�ks��k�ߏ�⇻w����՘�T"�2WU��E����>-X��U��#"�,���V�#I�s�֭�a��a��i7����{fS�����Xh+��YFj�c�����/N߼<+�U�q�v�9Gx�04�쓼ܶC$qZ����4�t��)=���K���d:��}h%C��D��"}�Z�jV�����7g�<������әQ20eەί�>M�
27Ø��S�Q�d�lm�e	��{�Ǟ�S�ٜW_M�x�&U�&͕P-��!v�1��������'��G��O~��ݴ`,1
"I�Ӽ����v�dICi&�W^{���y��-�3r����ˋ�h&��U���;������<�.s4$�E�6��V$38��&,;H�-;���nY�qx��W����c*m�6V�Cn������َ��3~��_p~v�_o[f/��R����7��3�ԛ�f�D�C�;2��0b2��Q��!Y��� 6ptpȭ��̪��Wl6��I0b��XWR�,c"b<�j�!�b��eP��@Ҧ
C��T�#F�Ce$i+H,_���OÒ��jp�R�͘Aʰ6���6�S���ϧ��H���UZ�an�(����,i����ޭ��}�Âl��]H����9��1�M���s��}�3WV?��j]o]���~�)�g��wc�e�4*1�h�1��3k�ۨwZ��{��_�p�gf�����hL��Sj����^�MӠ>��ʲd�~��>�p6go��|���zk�x��#�:U����,�ެp�1�͈1�^��҃�ݔ\�BׯО��>㺆��k^�<wטy�V�<�����B�X�9�DljJ�2�y,�L}Ù�od�{ʪN#ik"\��DIiЈ����#��y��_9���#�ք����xd� 2�,2�5��%�cR��*���
4Kj[��� F|���[U!z�{�n�<���)~IYVW�EU�����w�Ƿ?�.�=���!?��O؄��ށ1U`�ʣw�1Ơ��YVp||��߾�뷎�Y^����?�A���31���f�7�88�KQkh�5{{{��-`0����O_	���`��㙼6-]<�����Yl����T`209yQ1�/8:�A����K)C1�9NZ[�1�2�~��F�f����g�c��g��,K�WԤ�cR��G�:^{�6��6�2G}@���K��ϓ$A��`�l$�8ź��<#/�5b�S�p�!���8���.
�ce��@�T�g�3�I�D�m�_�}�����W�����9�з̆������p.v37]wu�we?/Z�D�f.B?[I�碑е��,pրFnݼ��w���?;�</b�7���<+.���y>�WD1)�u�*6��uB��j>�z����~��G�_����S�}��_Z�;��9��yL���*2e�B�EA���w>��g%Gܺ�*��=���'�z�`j�P��{2��f��ގ���)=�|[�iD��1q���a��z� �E��)�ڦ@�x�=U%hD4�5�c�!�b^�bi�@���S{~�����Ę������׵!�������H�޸��������|�Wy�W�厧�����SX�3c뼘ͩf�"��e���2�8��r!�����im�y��_��[oP�
�6E�#H�>�׾hj_�GVV��TA<�ރ�ϷI4.�����⌣A>4�`]�S�%CUU,��KU1�3c�;��#J�6	��	�L� ���n6��c@���i6}���N�Pb��,m�+��;`V-�=m�4��u�Czw�L���8���F ���;䭷�Ҭ7|��4�ŇTt���8KQ��y�M���c���w��tmMY��Oy���V!.�J��,��&O����� ���#����QM�Z2l�0���P{�1p�����'�!�[�J[w�.��ldq��	�b	l��u`����|���5���W3�sS��i��U�Q|��/$�ug�hL�O5��O��{����(J�>9����N"q�}���Rڶ+˂�m��*xpV��hEPcqA� z;�����޽{'������~?�^�;==��i��<�L>#��W���1B�v���WF�$Z��#F�,fs||��|k3���X��\��|۷�I��C4U�%����*��]�]�qE,<a��c�^��{��o�
1�?ϓ�~(��7=Cd9���c��4�k��{���zI��&��F}[0��l^���&�9v?{�}���u� m�P�2I2v6��+\��Bf�TH$��9��R���$��,�c��;;�Ȅ�}�I�4-}FDȜŕe�X^\�֎�y2c���׷vm �P7�:��i���^�l6�(g�9#Ĉ5��o$��R��c:�^�8�,-�A���l:V�����-j��.x��"Y��Kתźl�oEl���4]ϔJ�K�~��1X1��IŚQ��|>6Mͦ	�Ͱ�@q��s7�����X���a�v��2��u����6
Yf�Ǽ��?���&�����%�M�k���Y-*���'|p�ۼr��1p��)���'����E��Nט�U��������v~���-��AŌڻ��h���m�R!��AcD#��Ohj75��B8�����j*n�IB�y�Wc���p���|
��ސ�麧����;D綝�ɑ�|�"�?;�Pb�Ȝasy�_���G�7o�8C[��O��������N��������w�<#s.�E�v!h�]�{�������㏟��~��ٟ��E#iܻw� ��?�?�P>��c�������R���q��I>:?��~���� �/��\������E���B��������ƍ�_{�;?ߗ��;NN��ƍ�z��}�}�������_�p��R88�{ĠbrUo��S���~t��òX�s�֫���u���s���G�D�z�O7�u��m�1��c?}nL�M������غ�z��������f��1P_��m��v|���lk����r�Z9]N���q"�5�ױ|��^t�v� ]��aHJ�^��	�5l\�!%�:�b�A7��Z�:v��k[T��4S=D�]���[Oȁ����{{{l6���3�,U��Q
8�]G�帬��H^�1���vKM���c-N����e�R E�M��,O��ITn�>X'���B$e� �Q�|ĊR��]�s�u	$���u��� z�w��	���kD$�����W:�ڵ��*�����t���mi�T�Q!
�W�=�x�=n��:o��O��qvvA�S�y�8�q�͛798z�7}Т|��O���gV���S�������MA�1�	���	D���TE�r2�0*D�
E�p/FM*��I)��Q�@��ԛ1�}��v��'#�&�gX�oȜܘ+ݛ�s�nM��� yW߷�^H
����7�րj�5�]S�b3�t�D�Ռ�����?���5~����������A_#OO��޸s��52�ϥ,�.��m�Vź��Z��e�H�T���_���|��;w�5 GG���%��������Ł�ϗ�$�I��O�	K�b�ң?�|_��������E��sa>`���ê�ͦ{s}e[�u�C��N���θ�+�r��23ޠ�>�O`��6\�����{pq�^�*��9�rpq�7n��­��m<�߿������߿��Yy ���9?7{'{�4M8�}*s���b������st�h���ߗ۷o�p~��G?x�Jl��[o������&ڼțu�:0b�*R�A:�����Z,�mZ.//q6�����.F888���z��7M}��Eu��l6ڶe�Zqzz:������*6�u]�V�Z����}��޴�j��}J��qΡ���r9�С�k Ä��y�f�T]Y�	��-��H9�HfӢ�uE�<��뚬�Fp0�G�3��E�,�g�u'�9��ֺ��m8n��� ��W`�"��U_}n�<�����()=��`�\ARu�b�@5�����:t��ia>�,g:�{M�]��D�#��o��2U�>@0`�M�L�R��:B�8���쒦IV2���N���l65y^��-�GĘ����C��7�u�|qH�>���:)��e�]�ڌ��QC@0.��L��օ@<1z��h�Z�XU%�YEa��B�ئgx�9��kW�hH�P�u-.�8#lV+�͚�zMD�7-�(P��@��*��Wdԝ��k��"v�h#1P��a}�V���xQ`T0y�KV-�z�Ū�����8���V
VB�$��ggm����5?����w���y��1mW��6MG״�9��l�ӧ?��<<�es�M�K�2����g3���8�.�H[7\�^p��w�N����999MծU�5>t=A�g5h)�=ڮ��"G������l�������Ӳ,�l6����u|���p��S��=��&۪]�����r�;��$]ښ�O��a=����2}l�Z�����m6���[�4��:}��|�T�b�mNOOx��o��W<�����=��������w�ʃ!{!���,�fM�̾��o�o�w'�?^���*Y�AbUZT���ܓN    IDATET�?tm�'���J�� Wu�ie�Xi��^D��5�w$�pb���ցD�x%8a>3�M��=Ʊ11ΈTs77̚�n�K�����;(Ķ��B̬�U~�l����n�cC�z1!�,����!�.j� ��<-��b\�}p�����y�ESA	������tvS�l�A��x�ez�7U�����N���6yfo��u�J��d�w�j���;�w�6y�m[h�7Z���E��f�eM����ʽPU��.+�B���W�;_����(��Vwſ���한��o�f�ݸ1��ixp||���������Kc��l6ݽ{�����NOO�\�5�+13Q�1b��ī��mT�n�,�x뭷p65Ä�&��׫x���(Hk�dbY�e��͆�O�r~~>�����:�Ŕ����S���޾)��g��1�u%�,��z��qS�X���)к�=F�>Ҵ-M���-Ӥ�k֯{q����n�~��b۔]�!b�	�5��8`zoH�5�0<����C_tS����`$1Y��a��5�-�RW��z�.��ζ�=�3�R��:V o{٦s�ި��*[L1DL��-$�kX�R�%M����#���p����� w۴ب��1U��3�;���,�łX���5��c��H:&�Ӵ.�)�j�6������pǤ�����g��M��)��W&y���i �@k��9���J�z�L-��J�U1�*M}��ܣk=?��g����|��R��s.�k���e�;ڮN�[��'�i�@����զtl"�b!�v��3��{�����3N>�9���}���;���Z��4�II�Ľ��>=y�_�Uj3���#.�c��̥-Cg��Q�˜�N�٩m��Bi�Ϝ�磌g�G'��4S��2�~��0�ͮ��kԍ7&U�Pׁ��u�<1�ܹ���G�����p��W8><B�ao��#O�HF��C����7����ˋ�VL�>е��T�C���\_���FI��Z�T$X�b�zb�eTD�Q%�kC1S�̚��D9��Β�J4)�*JĘ`����FUEĨ Q�	���V���ŒN�Һ�v��-&�L碪��r�ƺ`:�Y/�b�[G�FuAr��G�k�����R�h�4�t��D5��U�#&s���-vf6�"��"��\��3�f%q�\js�l�XjŬ�ܬ��;���K�ɨ8��1뎉�Hې�m^��q��q����v�7Y�B6��n6�ʲ�ks���b����7�g	٧]�uw��]��?�*��]��<W�$�6"#:rwӃ UUq���͹�\�&�ҋr��k����w���ZR����#...Fo��b��dL9�7Ֆ�����5ɼ2�N�=}�5�E�S6lH��_��_:��	�h�f#z�u�l6�Q�͚��s�����A#/��Tӹ�n��z�x ��(1M�:}��@H���\0k2��r��T[1�X�V���چ��X�X�8��t�2c,&�WR�)M�����B�5l�5���z�����'Ӱ��&{
��k��V��#Mo�������.��q����u8vb���4��L�"�u]ӵ5]S#�2G�;p=X	0wm_���
%*u����1X㈴ĘLq�
��i��8����₋�%��IkȺN�M�\"m[�&IF�u��S�r��[��g��k׬�K��a>K=�����Ԡ�>��Y�DB�@$������'_�����OL�5�\h�!lVAl9y���}�)Nj?������4�ҵB��@S�ԜG�rۉ�a�gg�|��߰٬x������O�tWto�����K=�-�؂:�I��ᗟӬ>�C]o�(�!y�7��#��LA�.H���yN����֚�|9�A�<�4ד)�{�� ���Sa���bI�<�ٌ�|��w���W_���^����6o��M����t1����l./8]y$*^��(���-2�yF"^���ω!��~�]����Uc�D��s�XH�D4@��QIii,�2�Ё�9�s�:^��X�V$��#U'`�%s���	䑪�m�UM�լJ��mG��/ۋ�.R��9��2�>7��Ġ��� �b{�U�:���;�մb��"�;�D�v�� �X���"�Y��Y�c]+F�j�1��m���a���F�"�=�EQ������i��sYQ,�z����ڍ*j�|]�<���_�9���e�֘�]ˋ%p�������������;�A_]ty��&hʠ��QTt��KF���IÓeI����X�ض�JFY�dY�GMI�W�%���G������<�5OUU�v5]׍�@�U�p|]yMY���8�U6oMi�i���Y���+����O�!�9��#��������M[P��<=;e�� �E��s`��:`�_"38v��A�b�^W$ld��WٶOz�4���ټ�xHYY�
�b�Tx;��I>���ϱB�z.�Ki��f�j���ҵ`���5l��?���c
=E,Q=b�X6�ߦ����H�3=XN��u�_�4�햳X�<�E�
_Hդ��(�Wk1
��X:�(�,+Fˌ�����O~�ӧOi}�f�b��LT�L,y,yQ�9*�xYg&Q]Had��������euq�/?��Y��3�g�,�5�I�~���)0��)_��>?��g|��_�o�;X̚�fɬܣ��j��_�C��/~�j�%_��m�@�`G�/"��Y��1F�&�8C�����˧���D����%��4W�A�8��2�|�!�D�"��߰<�P��9O�dY��U��!ec��~���y�� ՙv����{�n��c�_�6c�7����fX���dY/������o��ݻwy��w���;ܺu��2+J=z�f����������U���3�\�XV��lV�Xra��QCX��^���������Z??F�у���A�#��p�$1���hLMf2p��b���Q�_�W��!QP�H��QM^���9Y��ۜu�f�L��b����d�y�'K&�I.b2�JW���^ٴB0�"�)�N~��)�C�tmMYU�Z����QU3k��]�*s�͜u��1#��ط��?~}�f0ԛU�%d�r�]�|��c�Y��ږ�Q��W�f�Uf�jU����5��6���lfT�s�޽���/�l�ݻ�߻w�u Gu�LUz+f%BkĄ�D��$]�GP�\^^0��{V.5Zo�^�=UU�h�.�T�1z�>=���?�����o�4h�|�Z�z�M��=O�4�cl��vZmE��=�wB�� �nzy:AL��>��%Q���j�����jE�n�,/Y�V	��X|M`�<�7�+���2��1���ܚ
�5J�"5�u�=����!ڱ'��@4[K"�B�'�hVL��B������:�e;QJ��뼠�r2�h75�J�:b�p`ˎ�L���mQ0���勉�7��q���l��2�U�@LbOڶ��Ռ�#�����T�ٵ=�*F;Mc�j��ɖ4y��r��|�.�s��N��g?��䄳�?9�r�ĺ2u����9\��l�TC�^D�C_v�7ہ*����C>���'>C��e)����zY#d�u�1zbH�e-g��V,O��~Uc�ʉ�MK׮Yy��?��_��9G�ѐz��%EL�O�4�}
�<�F��<!��q���"��!u�5	XxLH�%F�@�,�-�� �ΧjQ��Q�1���t����3�������삾�rw��s�f��;�i1�n5���0v�߰�4M3j\��eYr���ַ�Ň~ȝ;wx������S�5'''<y��#'''<}�$IDbd^Udα��鹱�!����S��l"\��Ҵ�����s�ME����h�@HO�Q����'�*4>��:��#t�x�Z�HD4�&U���b�E�o���65��3��_�w�@V�bFUT	M��3��g�+	VEQfe���-���(������6_����w��	IA��-�K�f���]��B�AIsL�<Yn������9(ɒ�,
��84up�\��ǒi}�P_�Y���(1!�����ˈF���,��6�1�%��T�o����;u~����'����2zF��1ƫ�
	�mu�� �Ba-��E�et]Cy���z��Wcx���O?��Ǐ���P�8�A�T��\1J��tW�)?l�Tp;�wx}�����@�n:z؎�x�뇱��M�1�"�	1|�5��6��כ���r�Rt�b~I�;�M������a���6���k$�)�#^=�E�<g���J�M���\����V��CϘ��9g6�(���,Y.�����L[��:�+d�$1}V�zk�:�˔��6�Ib�D��A�4(W��q��A%bI��vQSM�Rg�������ᕛ7�_�Y��ҮVtю۩�	�����٘��,x��|����x�����!�͆��'�כ��i+��a��rA��1h20F�$]c:{d ���EAS.�fţ/�8y�����e�6�;3���C숱E	l��B!s�e��
�Ո˓UKpdF(r��j��X9g1��3L��&}3@DL�'�TS��JJ�9k�3A�@7�ov� A����JJGG�(iaF�,�e��Yb@b?���oۧx��9�g
�^~��n����fC����9oÜ;�����zF^7���a�If�u�W^�|�=n߾͍7!����>}������
>65��2��b��mq.�陼���e�q�&����1a�*��Ҳ}\z���ɶ
��t�-��ߢ��]��X	��q�$�g]�X�㚀!1���^�Q0�.��M�vE�>I>���l���׈��9�y�&��1cG�$ˠ���R�r���ɈJ u��yF�2��T�%�,f9�2cP�X�O��h�(+9�
K�}_f���l��|�N�1l��HJ�u�
E1��m!���9B�9���w�m �#��*���f�[%Rh�)�[���Kg�����7��w�����Y��k���άx�������N����������0ܼy8���g�<�mkNN������/��p���[am�6W�����s.//��`)B�� �)?ܘ�"��=�vR�C�7����ԎcwB�J��w������x�i/d_��,i�+��~ۺ��/;�=��{�{~�GR3���<�Ry�[6��V�`�6�O5�@:z4
y^��w�|V���M��-Ѥ~��& 7'C0Q�%7n�^�7nQO�<%����21��~���p�$M�V��h�5�Ѻ������,�Y�\'����C:�,
n�����Y-988�ެ҄�@�Oo�Q�$�#�{�=�~���{ұ����$�1E(-i1r����ʶ�r�?��'Sˏ���muM�u�[%�k�h�v�#OA`�2fW�$��X�HP:�P:a��G�u��k\!�'Ѡ�2wX�<��AN�Z�]�cj1�ơ:y+�u��H,t��(���Pa�$pb��A;\JBh�cRP#�}�qH3�y_̐�}^���~�+�kwG�7���u=ʑRox3�q�5e����7��{wg~懁�\����|�[��7��1��'D���3�e7�u?7m�]�B�D��XI�<�Ec�n��J���Df�\N�k����{'�="�:��ύq���e����Σ$#�:4B<6sxBj� 6��GZߑ�> �B*�I�#Ĉȝ�� �@��f�X!w�Xd�e�0E�Yr�a3�3��f1��t\� A!*]���:�}�5����.�t͊ns��| Đ�m�~���@^D���C�v[>��������:L�UU5� ���p�Х�S�3�/f][w��NC좏A�uU+մ���<��o�7��o���%��+������8���w��l��d��[�$˲dnC@Fd���h�Q!�4��Z@��4�Y�H��;�l+��lQdS$��*��>��{�W�����[,6�d�[\��{��s����������:3Ea����+��V��pe��$�*���6M�Ǫ�B)��#rt�<R�nx��>[�=���bI�?����G���`�e2�\.Y,}szk-��m���1m۲X��*�d��n���tQ�"���X�'ɓ���ٳ���/=�OS[j����%�"*>�inO�7��8��V+�QFf�$����c�Y s������{�?�'龒/��M��E�/]�D�:}�8�X.�ƚ⌣����^~�+7o��(�{�n'G4�5���ڹҝ�q��2v�PQ���y����-�w�,�K����R�J�㒋/b� >��3��T��v��Z�b4�=s��M^}�U�I�T5�Uloo�2��H�Ef�Hy*�1����-ٙVYgm :��m�7hi��[��� �!A"J֕�:E_T\��ʁ	ˣ9uh��꺽tr>�1�>t�!aRf���P!�+|�$��&֩O�Q�' ��������1:�I<Zi�*pc/v�`��v4�%t�U��6Fw�����E�c�>��
�g�&�;#$�EQ�sz�|��g{q|�kG���u��7"���+wS`$���Ʉ���hc*r��f�6@r ��>�9:����@T'	�x4�{߯��<���(ǔ�s�}��yR�Խ)�&b �،Q��I�Q��y/$"X�is
(��z�����fٴ�I�ת����K�M��p&�&t�=�x���m�#�Yg�T��x���!�5e�h��LG kM�mn�t�kޣ�f6_���Uv>�;�+�R��&9�J@ɺ�(ݣDq�����z��=)8(�(�Qh�O
o�|�4N���m��ku�g%)�b�7��v�g����y8���6�`�\n�j��R�a�VƳ
�� �ˣvw/���G�������oE��W��cV͌�?�1<�i�Q���NgGL�SƓ�
SJq��5���o1����8>>E)�1ާ���½C�^z�� O��4��S݀�<��M<M
k�|/����~�w�|MӰ���Ç��U��H�>Csr�À
��D���dZ��-"��c��e��e�x�����I(���ւ�&�Ef*xT�γQ&j�)>�B�&�:}�_�w��g`�g����*?EP�����Ũ1Z�)ѡ�Q84���*��U��u��	%,������� �#C�u=�t��&E>��[(�͕K/s��_���i�@�\���V�d-[eƃ�Q��'(}�>к���Ӵ�n	��V���r�EE^��$��'�a�jE�F��<�,6h2Q��튑��Tx�Ȳ��Qň���k�����OJ����]v������������#��=Gh�dh�O�=��l��K/p��7(��x�-��'ӆ��.��㼦�9:�,��� �
r��!U�nF�d��	8:�E ����ۼ~��ϗ^�1�VGp`u�!J�b�fg?���},�cE�� 0�.����%�	�Z,G�n
13��$lN���.�$	��1�����R"T�l^;�B��0�D����9�=�E)��!�t��Xaӱ]G<��iC�,�Z�3KE�6�M�~�a&�5m� �-�uEU�(��_���{ h�(�	�̡E�#}(pz�b:ً �$X����h�K��B8�+\]Q-��nUL9��<\���1h(��rdg]&J�>Z��fvtS��f��"���,�K�0:��y$�Fk���A��W��9�w=H.�H)Q�vx�����������c�AE
��cg��\W`��|ۯ��1d���sWW� �#m��s�(�ƪX���=H��#t�_�����t�������ޭy�!�u0�w bj��߭�Xkh3EU�m�〻@�n���
���g^��V>�˗������,����QZK�����/�M3k��f.�,��[���X���~[^{�TGs�:Q&[��G =�/^00R����]�ܹ�������l�����[oq��-����s����}�:y\GG3._�L��ܹs��x�o��o������1��ǜ��Fo�5�D�>�mvAaRl?������3Q��%�q�<�x��ώ�������A��/y�q�$ �g͆)���Ǒ�i��p�N$����˼��>���~��l��tL����nT�%�h¨�H��]���Q$ت!�    IDAT���ZK�t�g,΋&�s�
�����cn����I�$(��	�������C������w���s�Έw�����M�v\'7�g�$�j�(��4�(��mFcW�&�#U�f�e?�lΡ��t��j"1=�N/�E})���9�Ʉ�,��f(5�����⠦*ߴ�TŞ@�s�b,�E�&�u5M�hh�S�ȳ2�.���G�{��K��c��9�u����1%�^kF�6��!���v^��6� h��^�0�D�[���B����c!C�{T3�H}��#s�og���^i��A�1�����k͙�cHAm�ޟ��M_�Sy<�;�:Q�E1>�Q޸����sM���.�����m	N�:C�eUD��kc���7�o<J"�w�d�e$�v��܋�8�*ˊpp|�����w
�G �������?�C�]��޼Y��� �k��R��cVr�pV�>��5�����.�"G#4Պ�Ǐ����������Xr,QH#��R���n:����)z�"rC�B�*|�=o$i�����t�J���l
��0:8l�A��c�{��QA�<��8h�Fbi��l������,[�xz�*����rU�ZF�͛7��sz:��dƅ��Oڻ���uǁ�vc�w��^p.��<�êm�yG���?�����!��LS9J�H���ˎ�prr����v&ܼy������i�k[�	�CL���E�<����� ���#tabׇS8��Q�t\��6�{?c�o��yLrf<�����>�eY��|��QJWN�v`����D��<��g�1�Z6t��-�SB�ڵ����"h����ƍ�@�bQ�B��Oiac����u�u������i\gl�G0�5=�xPg�ADȳ���E�����Qx\��u:��Е�F]>m#�/�QVG�<4�9B8+~�;�f�A*���,������"Q= �MA�������ߪ;��<�FY��:��˝t��$f�b1�CY���F���mQ�>q͆�2+#�,�."�u�w��Y�ʺk�#73�U2B�m�Z�"�����o���j9�EaQ"���m���ҕ�!�6C@+����޵�Z���K�$�E�G�j�/!:h�1�`D�&`\��YU.\����;w�0��1�0�y��1"���1���K$�:����������'�'�y�7����aLy�/ے��CO�i���Mj=_�[�B���Ң:�H�{�����s�>R
$�u�Dzr������.z�7�{�5i}���{�|>����u�L��P!`MI�QAp��l	jF�j�Ν:�<~����ׂ��3.�paY���`�ym��\���s^ʳ�~wi-�c�����e���)M2.^��d2��e��:FZ��!�����f\F3���� &C�"+�vDլhR�����I�����>[�-�Zk泓/|�Cg9��ZF��ɄK�.���)B���w������D~ga��$�`�eU5� l��q��M�]��x<a:��X,9::���������+ ��M�^���3PQ4f��<���Ǒ�qڲ�k�ީ )5��1�'���(���҈�B'���X|P��<%����FcTWr���+�Gi�o�t����Q�%η��b�Z|PH��wxӤ1K �.E��&�4!X�b�������L��@b��&�,�z]�s:�E�.j9�?e�"�v8w�E����z݂5����G먣���UyL�g�}�I��EiqU̈�m��AME����V��Ѹ�W�9�ۣ�3�#�[��w^x�;��*S��sJ렻�k:r+
��'���{�6Mӟ��Ǐ{��h4:3�����t:�,�� \��q��3@+=\=PROO�~�J�{I�A�.���K��	`(�YeY��ks�9�=˪�"�@�QJ�R%�D>�ha]������'���&�,��$��v�������>�d�A9������~x�ӓ9[�����Q�)G6��E�ꆦ�c�$z���wTZ�z�ꊐ�wݤ"=Y��l(O�"���2��ֺײL �L�4��	=�{>�s������^�ҥKL&��S7B�:ڦ�Y�>�>�t���kb�m{{mjZ�ԡAw"��r��k���5�yub~�l���X�go�y����km ���ŋdY���Q/���Q�����Y�ك���O ̘��vQ�ƹ��Zr��n�x������3�{~kh[χw�X�8::���CNO�q.tѯQ&��:��d�h�Y�#%��E�b�61���T�[�4�o%��p(/��^TҴ�V�d�H�Ġ�{A;���(c��|���V�C��DmE�AD)�h|z)�D;�Ĉ��:u唏Jv�p��w������N��|'����	^�(�g��A�V���V.x	�uo&j�k��@�j� �R38F%�{q1L�<*"U!T�~QJ�6fuナ\� ��AwaU �e��Z�R!�(o��D�;g���5�5���7�m�Ci�^���~,"�d��cT�#c�_TҾ$J��.���D����+�>��ݰ���p73jn0�AS*��.�b�\�΍�e�|���I��h�?$�D�;���ӓ������dIѮaĦ���q�@�{�8�É,�8�ӳD`��ϥ�0�Coq��U^c�!S�p��'-|�&���`C��� D�D��mt6Fk������H]��{;���(�mmAS�hcQ6G)��9Y�DӇ��w'��gr����y�g�)�ϸ�O�cl3
� +��5�c��tM]S�Z��>����6#�
�wH먛��ZRU9M�p��iA	YQ��w��tBF���
��h���D�6��	"���f�yk8&���:cl����(Pb�nR�T��g�\��ߟ�'���kU��7�=/��uv���F#�˚{��������x����rA�BuC��y�Q摧�"�Q�b������x\�}������4.���*���.�j)�̓+�U�#�#"!��˃3�6�B������Ҳ����T��SA\�ֵGG{˽�����RY�}���De�5~���Yf-#�m0bt�G^S*t���8��ʊ�hU(��X�j��)�&JFi�%'�$=�L����z�u�M�h%:+�P�X<+�m;�����E0
e�Z�VDƙ!H U)%�U�P"�(gă2h���H�2�J��A�ZKP��֡PblP%�5�eZk/F0FBQ0� ^,J�,ӡm�>��Z���Ѫ��ӣ��2V�8����Ց����Z[?�,܍�dr�v��}�Mu���Fo�컂:2YvA!c"�[3�6�\p�ek:��Gwh��o�@�4<~���>ƌ�q���0Ĩ�V�>���9�ٌ�ju�T~a8mxF�睴��lP���P�~pm����I��a��a$q��F16�_�K�mʒ������OZ��l�D�(��f$@G~L/S�����M�w���{����d��$[����f��ݝ��&v�(�y^c2�9��}�ш�h�<� ��{�6���Kkr�9�{Q1kL�oK�hkk��ׯ������#<xR��0x��������-�|�2�Q��|�ֆ�V������=:�{��p^��+{>��3M���%��-t�R���u�z�g���I��'������m&*���>^�o��;o�����!��
�'�:[W��6��&F)3Ma.\�!/3&[1[���y�_�4.��yh�Z{�B+�.�������v����+���b�ֈ4���MF;�V�΍��b]v�4�,���R�UVm��.��x5*���3����o���_��Q����O�(�~�w~'�����z���۷��۷�J��}�������t��6f��R�c�ƹ�Nm�k��f`�UJ����{�L0�k� w�X�TN�h�>�,�*����*��\#�l�:d@�dNkk�C�Pʪ�����D9���s6h��Z���8��1GΙ\i��֫;T�+��*��Q=��Tv$Y�a0fi�ʴ
�m_���AV%e����t��r)�nݺ%���8��Ng�ڪ9Ɋq�> �Qd���Ն�ka�X�e{{{����������wI�(�F��szz���J)f�Y�oW��x|��ؒ,�đ�`f(�.�O�g"��?M6��w�Xd��3�9�ߔ~;����6
9λ?�`/�ֺKu@���Q�1ژNGS�N���}�o��_W4�Q�Sc3��N2�����۟Rv�q6/�F�	�������g?�R��|Ч�O�*;����"`C�+��˶��ӊ<˹|�ba�Px����b�xd���ĭ�H�{)6gw��l;�T���k��
5��Q��싷D�I4X��"�T�2�s��Ms��x|����ŋH�O���$SJ��|��z<���ϕ+W����㣏�����hm�K���!f�(W�5ň�t�h4�����x�R��|�jYc����\�x���s�}ur|��T�Tm+�r~$J���EU��AB0^���ki���Z{�6M�hT��f��*��F���fbmc��Bp&��[���=���mk�x��znL���҅������ (
;�sY6��۳���ܵE]x_Ε�lQd�z��������ʭ�n�ɤ�>�����7.2�im������ڋo��}���X?��P���M��,�q�X\�U0�h�[��º���(-
_�F�bE1c\��s����H���Y�H�@��X�\ �i��~fA+������ked$^��z�DNuΞ�m�>
5��⼘V�4�B��ʚQ�C}\Uvvv�yؒ�upppr��α������p#��TL����0S� ̛Z�(T���;��{���_����QJz�w����ۿ�ۏ�.��o�b\������-�7�#����"3�l�o�V�u��+˲�%�#�u��UJQ�%�ժo�^�6=����CUU�C��]�Uz^�^� ��� �
+��<Ŵ�a��@Z�=��E��(h۶��=L��57'�=��x�5Z"6U��^��%���15J�v��Uk�8����F����f�~Y�(�δ�Icዖ�I��kK��g|��f�=e2��)�4� ����	tc� 7e���Q\�ckk�+W�2�-K	䅉�]%�/E�Z�p���^<�|��ޅ�4����qɲ]��~�yE����bу�ƹ56�<�_���ñ�RcQX:�#�����m-��˿��_������}�փ��gJ�G��:g��*>��ӣWؾfI�u�f�b{w��w�f�4��X�������ϊsǺ�?Q/"�0F$�#1p�6���~Y��}=+���:�_����ܴ�j�Y]�MK|��y9͛OK����,��y�h ��^�\�l�e9�aݖ1uu�	����Ɍ%���;�$x�ݽmnܼ����'�����&��"0�n�H�R�՝͉�c,Yf���t�r��������a6�ك�G,���nX>>���cw�?�^�tq�T�#4{2s�}\�֞�.���i''ƴ�͛�	ʨ�6�������o-���\X�.��_�z����)��śo�)Wo�R@�}��p��������խ[�$��?�?���۷��q[����i�[�n��&��81��G�p�_v��|{�j�]��6׏.�ӫ�h�ԓ�AƩ���q+���������cK/n���T`��v�%;ń-�VK���YQ�e�L���Q�y���*7�(9����ж���8�Zoy�m�*�B�h�5tЂ<��h�WZ�v��o��.m�z�o�����t>����Z!�F{��2�����R&��y{4�O��T���O�a���_[��{�;�V�daU�em��j�7�~���P�h��L_nr!��4;/�;�NY��ʟ���j�t�Y���9���
'''����^k:�TB~�bك'�؆*	;'�2�ȟeK��	Зe�d2������O��[C~Q�����$o�sBw�ӭ>*����(3�>���u��h�B���Og��Ιυ�����|o�"�/_�j>D��Gk���}Ї������/�&t��|}���-���:��p(C��2�d���|������obm�\����w?���lxZ����Z>�w����������E��@v�.����1&>G����Z��OKe�Ά��������$���s�k�d����!t����p!"�����8�
�>�E�;ֻ��x�y�w89��M�@u��Hj�f��s��e����L&�y.Jf���?�c�֎�jI�liZ��DJ��X���/�)F�����rn"A���eL���M�����?�c� Z�Y/9�o�������7���|����}�7��称$���R�����۷o���}��Pr��n�|�p��5�����0|�ߔݺõ�b�r�ܿ~]F���|�W���C��pl ���t���N�>��ӝS٫���Ω:9��s6|��U���?s������y��ξw橺}��o����<�Gʚ�b�]���՞Blh%7Zc�A�`}�&`��k�h��k�w�F<�����-`��rN$h��$�L5}R�i8qE��QL^�P�15�NQ������������2C��tLÔ���kj���gV�ՙj�/Þ��?��he�dfY�Ot_��=�6�
8[nm�F�hm�6�茠3�����ϫ���믿��䐏��ؠ� ig�OS�𐃇�88>b{k�";�\�|��/���Ǐ1&���*�;ϔRԝZ{��t�H|��<�w^Tf�K�u�M�(�J��/�"��k�dgg�����?�0�y/8�e@�v�w�i��"g{� �/���׏�墦i<u�X,*���"����Odϊ�mF�����?�g�<ǻ���p�ĭ�4B�]���o�7�����������|7�4�`�Z�4v��4k���QOK�k�d2�{��f38==U���qۺFIl���E����p:���	�R֒�F������iZ�����~0|_YgO�ގ��O�?z��I����g�������+���%s��<�ƨ�J�C����R)2�Q�Z�c��nMQ�aUk��eC;�K?�;ϔR]A�Y��M0��)B7�L��<�{^�d2��ݻ�W6L��xs�J�F���1G_��tނ�,��������%����Z�96���4�*��E�X������|�/���������گr��>����U�B�3���̎�m�v���1<~t�������`w�W.�@fe]l�w�OM)n�Ϳ���i`o�vFg��YG���d{o��f����~�G���9M�8�ɰy�V�K�>��ݻ��ҋ\�V���u7��d�b��,+O𚂍9dy�Y ~��=o�w����ڜS�c�,J۴0P*n{8o?������4�V+NNN��&���cҧ]�γ���
���CB�y���h΂�$ӚR�%�{i۶�C���'�h1����g(,J.�c�Wa�X�Z��d��3<R{q6�^�ܮ����m���৛��ʾ4{�]�������r��ҏ�׳�LByn��+q���J�]2�c�$�`:O{_Q� k�6�Ki�a�5�!P��_.����V+����,y��^���i�i�3�жѻLಪ�/�����yD��'"}S��z�I�y-ݯ3i�n<E'%�)�����C2��6.\�7�7�������_��`�b9c����g��aC�����֭��؞��۾��9��Q�m싊���o���y�/����`��˛�g�=sJAQ�i}�,snܸ��70�PN�������o�X,��#�#vDц�4e��ʐ����#>��C2{�����or��/]�i�?�׊�d�	J������m��l)�5���ߟi���cꪔ։��e���\9
|^��M��2<uS�C��4��?+�w68��{�ɘ��^P�X�����Ƭ���Y��3�ǣޑv��Ѩ�(��Չ��RH7g��hC�EY���2�2U(�[�!s^�9���+�[b�&n��xG�2[��X	�f�F��|�t�Z)b;�4 7���;�"d�҃�"�	��7�<ͳ�\7ӥ�{m��)�ato�In�tC,�3&�oP)�w	FiA�.    IDATӾ7�߰(%�y7���h;oR�=+���Y��t�S4�y�3��m�c)�O)E7���Y���7n����_g:���ጻ����!YfP��9(-X�	ƠuL�<z��*ߡ^�ܿ�|���'�FP%����;�?��7ql����.��9[�z#}��4M�`y��5~����|�"Vû?>������?��>~�̒)�hd�@��Sa�Ay�.�?�����-9x|��l�h4�,&�W(,Zٙ����7�=o�����p���,����9t��Na����f��y�O��l:��U��c�ٌ�ry&��|<��[k��f}�.�S�EQ�Y;����4���c�t�I<�bKw��'`��G~�24MMTԳ4�w>2A�w����n��~�\�W�sjO��۷o�����!�V��^�6<ԙ�����iM�7Z��(5&�Ch�p�I`( �1*6D�]oǓ���dO{�Ҥ��KO�WaO�o��H�Q�}��[)�Wo��䱹X�m�^O0���,��Eq���ާ�__��霡�7k�N��p.6d�&��O��^Rᣏ>���j5�YΩ��Ѹ@���V�k5�讗��Ǉ8_��c��X�>�YE���t�U��F����ؤ(el�A*�\t�3 �<�T��F��OkM[�k����h�[o�xp�.o��gܿ�6����N,�<뜥��tJ2Z�@k�.62OQ�?�˟��g<f�#��P�<'�3$(��i��r�i87�\W���6���������O�<?3G� @KmS=1ߧ�|E`������t�S6g<#"=��yl�����ޡX� �@p�.�F��J89>\GJ�fT���m��bբ�� �
�VC%
Oӈ4M�
�[�L�Q���vF�90����)����,ٹ�Q�])k3/.��Pg�}O���J�Q!`�����d�ė�b�C/FDX���Drvayz���8�D�6��":	�=�Xy����XP�0�����0�;�,�g�����E)�{iC�/Ҟ�>P6��I�NW�ŧZ&"]�óܸ4�b���µt�)�lmm���͏~�#�̀��oO�u�B�Z�� �Y����s���|q�X�W��bww�</�>�is*g�>��,�"{���oq�ٟz�r7>7�8&�	����~������7?�G�<E�S������kY�jl&��S�(�w���ȩ�#���ׯ_�������cr���?�B���3�u���
�}
�S)c��E�R}TjHU9�c�4J�$@5�N�N��-e�Ζ$��|>�[�����9�a�#�L�,���<U�9���L��s��i�_k���.�l����YUUvMJk����s����s����S���i����Yn�	M���Z��nf�}��>z�b���g��}������~5b�߹2��������B����4���]�[�Xm0��j�kO#^<"�F���-1�:*yV���U�j)�:�������kc����<�ŝ��j�a� .�u ��􈭭-��'��R�5Vk��8�Hal���m��2�=H�w����
)LqH^e�Mn���� ��7����0�>�i=�d!�I}}4J�j�r ��/h��>��� �8�ٚ쓛-�Q��&4\���G�,���;�2C9�?~Ŀ{��</��?<,
l�i١�u���/��ͪ�����7�������]>:XB�^�ԒǇf^�ƉB5�,���	�v�-7a��<^=�n�r˪
 ��Ni���g_�O�JYT�G.��R�j>CG�ۓ4C��j��j��
5���|�Ο>)�n����F��j9��Rж5Yn�ti�w����?�x睿���nG<<<��m#���B>�3���sC�t4M���1���$m<��=3(�S�Q��ի�2�@�C���D�z�jǣW-A��8��*�0�,���S�4ԋ9�լ�m
<��&�B�0
�P�סu���in��]�������傼(#y�	�B�`	m�$p��un\����.{��\��C�@�\��T�GǏx��!����v��Op��K�0s-��2�C�U%˓%EQ����o�̅+���,�(Ǹ���vI�.��ӓ����]��>��	�r�xOfGhM�'�ھ�Py=�k���<!�E��W>�Q����1��h�s�����a:����@�E��<��IAr(�����@C���-J �Q�f�aœ�����Jk��y��"u���N���Zw����P����xoG�z����Bi�l�������WK7�������O���~��\���o���=�2f>.���j��^cj����5֢۞ �4C~�Zb��^P	��k3D�D�C���Z�x�}�6ӌ�s���\��e�G6�|J�*�,�X,,f�u]������"ҡ� n� V���(Sqq={��@Қ�xn���m3f�%J��Ձ�N���E^���SLE����Ÿkf�Tt(��歚Nݿm[=���½{�x��8<<�Q�=��hU�V�cMp:>'*�d*�x|h#�V!v�t��QT֩<?;�ƒ�%Fg�ҢM��nɣ�����)A��Ϣ��o3M)�	����߽�|�[����V@��ҁb�T��}�"	���"Q�B�M4����{���(���X,���u��^`o\P��`��9_�3�/m�B\�t�Wn\���q+�ݿÝ��`��j(EfKP��n"�����y���y������&�g�2�h%T�mUst��;����ŝ�����4%(KnZ%,]|V��x'x߲XԼ�����_����Wٿ��YD7�x�i��+����f4.�t���O���(�5�J��by��<�j��ß��ݼW�"��66i=ß�s����q�7�g���3���y�X�VH:x%X��"�y�T"�{�ӗY�ʾT;�����w�w�R��j]XV�f�ng6�&
�ɛ8I�c����'GqR�s�s)-���#�=@���
��k#�>����,A{�Ɉ\�OJ����ސ��Ep�6�DHN���x�ŋ�����?11}��������*bH�D%@�z.�����M��"�i�g4)Ȋ��������A+E�6<>����9	
c�و<O|��H=��aZ�1���,�Պ���>"�:�y�5
�"�4�AO^(l�vEۮ�"A;R"@z�;x�"�@��1�"(�r���+��w9\T,jG��,��UZE�a���go�c�a�~W<�bXձ��6�ۮH�K�� �G�b�QxeQ0Oy�k/�5E� �N����� l��2���ɚ�y����y�+��/�2�ܼ��*��>b1?��g���2d��ʫ����_�����^���S�?z�S-�q���-m�	W.]�՗�ί�����.��۱���)Ah]C>�c4Q�w���^fz�
[��x�wx��~��f��[�LV /�g/�t��|�;|���foo����и��ű� �5�0��^�0#���������;�NN��PZ�q�i7u�L�9�)���?�o��͹<�p�t�a�es�ߔ��<��-��=�:쬳XA���������n�h��X�쩒���X���$��|��Ai��u���kk�1z�m�A�A	��Q8g�u�IWu�G)Aa	�j��;#��^��<'���R�^a�Le>˞
��0���,)ҧ�ꏡ(
F���詀��MЗ������C�}q�TmC�^^��#��.b
��e����%`��Y�,�Ե4��j���Y��������������hM�+DJ�(�#]a��6Ɠ���5M��iWx�PZ�Fx�vh1���6*�"|�Y�"���`���~�%����:�V��h�Q�z[(�� �Ƣ�b�d4B�15�X�Ed5>�h��]L�J�Պڭ�m�����h[b�a�j����7��˯p���fww7F�f�UL�F :-��ŗ`"IX{0?)�6�[��ï�������������d>;��Š�k�< ��1Fs�����7��.�v�l9c��Ĭ:F���-uAqq����_�W�W���+��&�^@p��r/�����/��7v(&Q�6*�����T�C���8/�G�ܸ����	W/\fog	-u�6��и�v9��
�������gS��0.�@��f'BL�~��Ր��C����E�Σ�9����S@�y������y�o�3�u��:�"H�v�!�J@9	�&�p��͚�~����?����o�=��1Yݢ�Jk�k�2c�dJ�1F4�#)��#h!�yDp.����ćF��Ak,��`i��0x�o�x � 7�~'��>�ڞ�4]c	Lӿ�ņ�J��$�Vp���{�r���Çgdl6���P�ŚD����F�I�9��9Z�Bق����Q�y���Kr���LIKp��b^��(���2��5���D�5dV����P�U{���J)���L�#7��ޔk�.q��.���|M�V�m�-YG��#�炀����F��4��1P�kF�l��/q�i�Nv8||����U�����,Fi�����(�mc�⪉�������zE�j2cMs�<��CPh�c���=Ⅻ�^����J��y��&���Q)eh�Z#�}����X�<�(A�`�G�B���/���OQ�(�c����X���~�ݷ��|4���m(Fc�|L�!
��,˹v�*�x������%���K<ZTg���%�k9��|7���)�\�V���3޽JZ�|t�YՐ#P9�5��������^~�reP
��������G�G�mC����/39�Ɉݝ�}��Qd}��J��ɊŲ��ʀB�|����v�{Ӝ�Y��>;�^�y�\<�T?�ZO��͵j��u����ӂɩ\��UW葧�� J�	��ҥ����9���SA�t��
?E�Z+'(U�km�3�kl0J�lv&2`�A$j�:�����K�$Yz����9����wuW?���ְ���%��� �=;o	A� -�!�` pe�2�YX^p�	�m@/J�!��GwOO�����Uu�73#��yq�䍛uoU7��d��
�73#22"�9�������-�@���:�Օ�1�Cx���Y��QL�~Ƹ~��#-k1N��_�����Q�ũ��l�<����9�#��:��?�������C'����#b�H�KPK9�������X.��)�E�`)�
c�we��'%��s��rs��Qb����I��.m�0�l0T�0��h4�Kk˽�q�˗np��y��g����7�d���_]�J>����EL����I�=J}qcs��|�p�ڳ)�8D��'�]���gOJY���ރF�g�J�i�PVfU�j�X�P�:b0����U�=��te��J��bZ����3 �g�N_�S�&0m��\�h4��2�3JYV�;����7���J�RVc�rD�=��PE1��¸������3����u~�������rI�l�}�}>���N7א���a
�_�t�+W�����-`�\����K�ˇL���/�����+��ʷ��[��)�o}��������98�vc���/"EQ�������y���v��8��mv/^e����]���"�)}�qWb���K�
ﮏ�}w���y��������z�����ѩ�ߕ�;zdH6W�"bQUU4�Z5z4n(ԟ����s�ν؛��Z/��}a��3co�m�s�)�(��9��t��J���w6 5mk��E�D�K���H�1�`�0,+$*N�%��@�Ā3��Y�!>d��Ͼ���\w�㶼�<��C�GGG�t�<�f0�߶���&�Riׁ��`��m���FM�%�sn�s�����J�}�l�Mݲ���ݻ{�
;��xV�.]۬�	+Ч��iq ���KBlq�d<�Q8<�5���8�M�֭�%.^��d���&��$�C�E�jf��>�I��"R�c&�{�
�VL6�lo]F�"QY��n�,����QU
SR�I���RU����!��h �jD
���\��<>�2������������Z�����M|���>{g��I"Q��;��u��-��Q��5X�OKA�C%�
'a����}��6��!"W�6D"1%�p��3�ʯ�:������K������O�џ�	��G?���vl2�.js��5�?�W�^��SOq��5F�1bK6����"BԂKW��ܳ/R�D,�ٌ�{w���ko������-���&��5%�bI]�4���hƅ;�%˺�	��{b:���~�+s�	� ���t�����C��}����,JN��o�m�����$2%͓�gy���Ĭ�`�QUkQ���drG���>�_��{,�Ȅ8�ʌ���ZS8k�%���%%�cde��5{����a�M�W��6���H�'�/UU�,ND�ˎ�Xc1ƥRf��x��]ξ�o?���[�,�lv�}ܶ����{�eh7��N���b��&r���K@&�ʔm�dB����q��1���|�!��S�o��{�S�<�g�c��˲�{���3k�K99��ǄV�u���>]�[#�2�&4M�F��h�h@KP�2������4��A����ѷ�2����D\$i�<�2�UИ��'��Պqs"��1eK�l_�m�$��u�\�b�2`d@�J�6�\
�p��*B<Fc�].8����s��]��T�b:	 ��sR:>��>9-9H�YV�)kN��m<��X�X�<�����&��J'k(�u]��[�˖��&/\��g^d���t:���f�C���Sn߾���>�����m�CX[P�wo}ć����6�x�%�ַ�|�
���8%�u��α�{���m���dv��{��[?{��{��G�!˦A���1��n�ܾ=���?z�g�~�ͭ��r���f�(+�i��|U�	���?uz{l]߼9{��b�:&�,�^�`���w���=�x�DE>���:8@0ƢQ��v��_E�R%�D���Ύ���~�'�Ϩ����vt8�gM�=k�;�^i0Rc�#"FL)��J͔eM�4+M�b�|DGa�Ŵ�8����""�(J.^�e2���ܺu���^R/	D���c�i�"��!�&su��pѯ�����2�=a��\[��s���#�1������ں�p������:)+&Q����س���0'GN'z�y�
���������h�ӕV�@J����ضH(\b����рyL�\)��M��[�a8�����'+��n��8�1 ��;e�Z8V�C
/+Mwo��Ꚏ*�7K��1�+�i*�7M�~�l6��n�[�PR/�(�sx�4MK���ǶAU���D�+���9��7_��o0�G�.��쀪�N��|�g�í�e*�ý�/�u��da����Cvv�S��b��(-�G<x�[4�&��WQ-9>�r���y�m�}�����K	56շ���CmQ0�����9�� �:A}��e�6*M�1�g�)lnm�s%��m��j�]��E�@?����@z��j��E�z�iA��2ٚ�c
��A5�i<�3�^��_�����[�mˤ2�P�Ĕ�g$`բ&�1P����s|��k׮��������p<_b���X�h��b�p��.�i����7�:GӇ��nP7��2�r�bI�m�lǷs>����xT[�-U��	��<9RSũ1W$�D/�G��yj�����y��7����!���:����>˷n�����~�мȄ����,%��x�����}k�rs|h՘I�X�{�������O��l��v.�{8(Km��
�p��ڐqU�Y�$�u֡eI)d��]�<�U��2Q��M�\��G+�(J��91����
��|�lv���>�	�BI�xM{��D��:\�J��9]�w2��t�MӜ���癥˝438ι�d��Nw�0s�n���}��u&��?���w>��x��d��Y���b[\QUɠ5qUFsU8Z��)��{̎7G���e6�i�}�w�������Z���Cb�b��Sɶ���~�V�6��9�H)�v ��K��=    IDAT�󂢌-U%XI�/�7��t������;<|pH�R�$6Ɉ�J7}:���Jr��pq4>�w���$�����`�h4�(�����Ո�0��T�w~���D۶�*�*��?{t�\��loo2W��o�펊���/��4�n��0;f6;b1��6e:we���;I��E�^(�c��=	��i�R�PI�
Ԓ3�U�O�7�O$QM�1��TU���:��,.��Р0�D�cQ�?#VI K��t��3��z�J
=��!�HE.	��ǧ�j�d�N���X�Q<�E4�8�H�^Z�5�%kEmm�$��j����t���ھ.�_1���]_4��4��c�z������L�X��;�(0��e2�P���EY��D�BB�T�W�bF�������k�w�F0��11��Q�D���F�Z�4���UgQ$�rY�U�ӦiXV	��m �S�0�k;R�i��׾��?���O:}���aDR1�ު(w³(�b�Aۦ�;;;lmmqtt�b�X�Ķm;�x����\E�{��Y?��V�
�e&�_�h�#��We��t~}��1�����1�q:��y���E7����ĉ��9�>������m�z�`9;bw{�A����s����{g���;;h���뀿[M^Ʉ|�Y���xc�y�Z�A���Bo`���r�<-���$c0�uK��>;:���!���L�3�`�vL4�95!�Y[1)�0� Q�<�xz��9�-0Q-�VT� ���E\ǔ��I�o�G~ͷ'���S�J6|��U)DS�w�UG���,t�p�V��(	�&�G�g"_�nO@�k�K�jQ,F\yS���ֽd��<݌@V��dEJt�
bH�;yIo
�����&�Fl�RFULt��$�M獧���g�@��1QM��Jʚκ�cҼ��P�t�"���,M���,@S���M ���q���5ޮGU��Ԭ�^`92c�5��n~����������"�ۧ���{#Glr���QըF뽯���u�ʐ��Ȣ��E�	��_��{���l��h��kj��%�+�����v,e-�25�%�cM��5���q�Ĺ%m�2_$/�A5�m��a8�
A5p�������H
��h�Ƞ�VN�3Eߟt�d�Y3`i����]nܸ����*���F���E~����_~���x�^Ɯ�M��h֍���5?i�R=�˸��g���iO�%j0�+�6��xk~ĝ�c2�ę��#�z��E�.��{{ܽ}���}Ignӵm�l��9W��k��m0�~N�6m۲\���6)S]�ǇH��mX֋�6��i��b!�[�,ʑ�M�H�,��(�/+�(!%�4
�8*�E:%z��6�3��$4���,yf�������мc<M޳�kڦI��8��J�� �rzA#^#�J���q�"Z̟�v�IF}��tL�t�F��
���n��u��Xm�+!�)�!/Z,��t/�x��K<��M�Ĕ++練}W��9���Mn�!��_����
�I�e@L�J$6(.�-&� �&�W:��*B�#`L��e��"]Vsx����[N���n��[�������ϓ���s]β��gK����)���0�/�1X�Iy�Q���c�Z��n��E�|�>f{|��L#VU��Ԃ4U�/A*��t2J�Z�B0�	>�"cbǊxr�+�sFՈ�p���)ꔭ�Lg�<����w���/pt����{��ݻO��:��N�/�Ϭ^�~�Y�,��B飣���N2�����ѩ��l���������s������ڧ~�3y"�p8d�X��˙A:I��x�ܕ��E��ΘNۗ�K!�\*ki5�8>`~t�C[a)� �6+0mM��ђ��Bʮ�!���٧��������LA�����m�jB\"&�
�u��䶟����Ҙ�#c�M���q�BL���R�T��K����4�,��X�5.U=),QS�L2>VK
�8Q:�����
N��Oq��º�C3�C����FYU����X��;�I��<�:�b�ˠ����}��
	jL-&`5M���N�������8�>�n��A�²��&+�&�E�H�`<I���\�P�3�M,�1մ��k�twh'l�E�I�ӗڸB��x���S�IxS�t����(�2(v�7џofVK�'KD냾�����Y������������r��Fl��}F����''�ϸn������*Re��,�ъ��x�4"̌m� �ۋ/BVߗ�c�'0}����j�O6�F�xYSv���F�R�
c|xR6�����e�hV����;;;���k��|�����&�	ՠd>����z�rѰ�l�8�V�&`U�,��Z,+�g�a>�����b���J��[���j 'U�4�c�`-gg@����,DO��;k@�"��~[�5��1i�������&�D�3����%�8l!�o!�
�@�HL��F�h1��L�E�4I�^�hh�TǖΔW*��^*�
E�S�$��İ�N����Θ��Y���ghi�b���,�N.�ze(��I�H,F�Nq�{�*u8Xy��{?�IY�Ic�!z��4�jK@ X�8���s1�b
�kH��D�X��[@�O��c�u�}&��l�2}��AC�}]���L{��r
�����jNd�;��a�3U�0E2�&U��@$1	$ÞH4i�ŷ�U�FD�">���b,���B��+�gH���;�]�ݑ���%1��0�C����I�Zs��Op��Aߺ�V��y��o��|ǘ��ׯǩk���~\����i�q���y��ַx*�3j���j�Xc�a�%\d��b���e�B�sA�tzE'�N��G�APO�����?��
VI�&�
]�\��c�cc#�lU���[o��o���\�t)�������������Y��(���T�N��*v<|�p�Y8Y�z�W���;d��3v�w�W�9�������'2g��Hh��h���Q����t��<��}���_����=�ɞ@m�]b�Jg!�2݌PR�Lh �� &`b��M�8am7%��b�w�o�k���_R�S
o�t��$�� I�
�J�4D�D�'��N�f|X"�슧��$���O�7&%�k*����Đ,[\WMG5%�� ��R=\���c�`�&�!�im���&��ݦ'T�vá!�F���\������`pj1e2ê�Đ�N�Q�m�����y��;o���k����U4'a���8�l]�Q���5�+�䟙A����S߰ޘ�?v�tw]��d�1�99^%%Y3�W�I [$+��eW
7{T��>g5,��[,�.�����9Gi�� �l� /�'����xw�+C,>+Ě�=u��`�ց�Y���y��B��\g,}g�c���+���`DUV8c�1VC�qv�"�p�h���wŪ�K���Q;�]�:��=E%���Ah�8#���t��-���v��y��:�`���dBU*GG3�ۻ�|�����Y,�Õ�i8��/r��e�����Ν;ܿ�}ˠ([f��t��2C���2c�����fh��B�n������g ��������=�!�b�l+�{�;�}ј>��][�+TU��]�P����6��EA-��o�-�2o�nM��dԢ>U��@��r5=�F��d�L
u:��&9ƈ+:v%�41R��#�׮�+�����	��~��VU�eC�6����/`�`]�(�.I:B��[ �`c��h}
����m��ʤ}5��>�QbL�/�`�+Ř&OԆб����;�I��bt���A'��+�>�?�yzb����*���#�rw������YgwO�k<m��+2�H�L�QQb�ћ�`�bR}��'�I���+ �IV+10'�;�poDc���KC�I��;O�|�������y5�巜��b��cy���g�}r<���g�_;+BsV�(��o}ΥJ5!x�5��c��	M�����7����:Ř�&�2)�������S���l��v.�����`&1�E0�F5�^�7���Ƙ�~���0��T3�<Bh}b%�j'�� t���hs��9f4����n�������&}t����՗~���[�xq����|���{�{ꕯ��dbT�|��+�NUW>Wg��+�]�;:���1��:r��#�����~ˬ�j2�uα������
�>n[���xU�7g��{�U��mR��xT<1Z����)�	��XpE ���`:;��E�	��]����g�V�ڝ�'�W�0�_�Aȓ�Y�K����d���pJ��Ԩ`I7�ѐ&�2�P#fD�w�ͥ-��UI��v�%b��u��<?�k�1��u����Y�_ak�E��t�DR �m�K�S���z�fxW�s���哄���bd�)7���@}�n��ۯT���-��6������^q��?IX���%v �v��4�$�r:�#���	gA�S�$�W�����L2���OK3�B�k��}���V�# �&��9,i0EEӂ1���@S3
���x��2��c��q3�2�7"C���K�_-�À-��Ō�[;4�R�kv'����fH45�)� Ô��˸�|��h�u����#��c��,��.N4�����$��˼�`��d��Ax�jk�p��.1�0��l�mB;$ĂڍY6J�~���­Ch:_)TlWkA�I�$1B�uZ�k��0� 堢�*|�Kf�}"�_�3g[٫/�Z��!�r�Hظ������]���ǝ
g$�B�S�Nk	�j
��q�H��4���E]����;\�t����������=�/�����s3�y�g����'�����v.���ى��)�߫�jEP�Jie���Z��:��F�;���3�-988�iF���!��>/�r���vvv)˂�tJ}����ի<���:�����c{{����GB�O
q�5�v,ow�����}��Y�3y^8W�;�ugc~��
f`��/g\gP�}���U�izN��az�?�cߏ=�!�I^��ʧ<���X
�)}�#�Y��[���Y�~���)���0L�9}?���HA�z
�Pز hK �k�C66��-8n����[���g,.\����|�%�ج@*�&�RT�;�`c�.�YR��;u����u�����\nQu�M=��=�/]WO���!ee�L�eX��;�0�K�zsG<s�;�Z�s/��rx��ͯ��W��
�+,�����~�[�7�~`o_��,��a�F8��J�X ����嫴m���{\�v��}����w|�W���Wee�����@#
[h1qf�x��ח���}����޸q#�m�y��"� RkJ���j	�Ɵ��q��t��2w^�	�3�p||̃���u�dr��G����?���o������.�����Y�7����ڒ�(�r�J�]FȜ���AOX�Eǯ���?p��?�K:��b�&�����	wbS��?z�EO�B�߳b8�4(<�~�-��-�b�2�z&�K�^�������|+u��3e�ѝ�~XىH*��=�V3]U��kҎN��S���i��o]�q�ϟ��ڢ#	�Y%���$��n�,V�,�Q���zl9fs��q���!���H���%֕X;���H`<��5�˲iPM����Г,�Q���%���P�����"4U�1����s�uU+X�5���Z���5��%�	��)�%A5���#�0/'�Q^�k�>%Jb���'2����_�>���l$��_�i�@-�������K����?]��ܿ9Y�w6Mr��
<>$������D,��ߥ������7�����d2����?���q|<�M��EӴeYVQ���HlU�i[��b{���e�B��f�n,74�&��H[�i)2G�RU[M��QU��VTN�T���:����ASČ�Ѫ�fs��e��px���k��s��U9fP�����N�ݻǝ;w�L&\�|y�ӛN��t�>K�;t������ߏ�v���e��������}��{���_�c��S@����ǲggl��j}���Q��S!���>}-c��O�2I�g��u��|҈����Gx���u���y��9�><���Re��>(����@��{��k���>���a�/:�%��D��/����S�K�� e�ŕ�np��5����̨�c���S�o]�JA3]2Y���_����M�B��*��O-z��uD1x�D
p�M�Z��hLY�ƭ�_�釣f��	3���@�E�Lb���'[1�k�@�!�-�Iv�j�	,j��骫��-�O�����\�u�����Z\���~��>@̥<�����=�#V�QJ�����ژ�)۵L��Q��)�[�<���/\��'���w�r6��?�F�F����g���x��F�>�H�=
?���ѧ+��e�\�sA���������E�:�u!%nȑ��*^U�*ASC:C�U�w\�L�ٳ.�RX̑+z�z2r��-<x���6��&��pLQ�)}�����u��i9��[o�|���z���:��g�2�9��Fn��C#9�7�����~bM^M�e���+�Ē��	[�uF\�7V�I��=������$�������r'ӌ����g9�kǄ���:)������}Z��^D#���]Z���Q}K[/y�͟���S�˘a�`p���ã��ܾ���87dkwL�i��-�������z�Kw��!������wߡnTO<��GZ�u#�@aS8�,u��:eoc@R&��l�O��1�_;C��5��B��s0E�+�P�T�ͤ�Wlh0aLԐ�=1Dծ�!����h��2�N��9ۍ��>�g��_�������Ҝ�ѷnY�w�y����Ǔc:�8{�����n�m�(+bT�&�o����ʵ�?�\�����H}�\��nx�޽�nw�b[��C���zUDE<Q�3eq��|��l�������_��M�֭[�+���\}�@����s( ��X�u��ߏ/����֭[���y����:��DD��?��qm�M�����j��F�eT���P��,����h��S�C�D-֔�XB�GC����������
�;W�پĻ�!����)}`��p8<�1�����H�|>˗�� �Y����ڼ�q���g���Z�h�rD�g�����w<-⪪��+�׿&�0��^*��=f)�(�~�TI��\������|�Ӯ��J�;���߫��||$�˓��'�\��˳&�_�w��67-Plʎ]},US����o�����h��k�|q¥���R�Qmy�����!�1�ł��+|����W����x�*�shU�\.�O?�?�ɏiB��
TQ">*MT�
;�nCD�g-Zv�%��Rv�*���m[�!/^d{{���ͭ{�C��� !�H*|]PT#�	�(Y�|hS�{R�$�HO;7�L&���7(˒�tʻ������^i���c_�@__j����c�ia݄߯�;�{�f�8��eM��,K~�6�ؓ��k�4�C~���L�\��'�p?�?8�z��O_ڽ�Еû�ãoq�������j��h�r����[���h�Ϭݼy�ܺu��n���op��ݹuK�_��@�y�62����U�P_���o~��͛E�M�`n޼�_}�U{�?������~n޼i�� ������z�Bw�N/\������E�p�:���������Z������GGGᥗ^
���w�<�����h���=�;1s�F�CsT�&����#�:�(�ӝiW1ã*X���\��y�7�/�گ��y���b�Ac�2/��-�����{R{�w��Px�wvFf���5g�<x�ߵ���qL�)���`���$\*g��_t��y+P�\.QMY���'��V�	����S���~���7��-�� ��#�r�9�ڱ)�I?`�Y1ۻf����2G_��2w>�
�/��ϻ�?��!��W{Xm�g����N��bwW�    IDAT4�����#�#�[�O1(6�r��(����;���䭷ޢY(UUp�+7��K�o��l����H��1}x��������oػ� �A ��5���BU�o_��Oږ��i��!��t��6b�ٚln������K/q��U�����kNk���h�����l��:L�lm]��s_g��s����ǀ�M,�I�ڳ'��W�~�:/����ܺ�Ç�<|��Tbŧm}��^�2��斫>��]x���ni���]���Z��p����e�z
�|�"O?�����)�W�v.����u��ۣ���xn6�Q�����L�b�+e��Ԉs�w6P�!L�o�����oKR0����s�)�[G
��`�;qoq���u�������9Y�	M�������^{I ^~�u��n��@���\}�+����Ķ�9޺  ��L���y� 	����tl�) �	5Ќ���rA�����a	j�_w�E#/����͛���~�e�������a�ؿ��! �H|(�O��ݺ��2ڑa�?*b�{��{�˲�"��Ht�;Ｃ�������Q�����*�(��XЗm[ԧ��"RG�V���q5	�����V�ie����{�:	�@c�唷�~���S��;���[��S��s1�#��h%�=ku��t<쭷?Zg��]}֭�ֿ���yL��1�u\^��_�X�����e��gn_{6g�>�=)@���p�դKD4yΉb���c"��H�!gN>��i&]b��~�_��3}�x@��:���{�G>z:�:�/�b�̧kc��ܹ��]�Ե�\�x��4lo�p�ZIQ9666Mvy��wU��o�5~�����+ϲ�<�ǲ�y�����������}���6�MR����Mb�)�Ոrc�_�֯����o���t�ҕUJ�e5dkk7��+��7 �@m����ä�>�|���]��$F��f1]�8^��������o�w�"|���⒢H �(
&�	���\�t�o��5~�~�?��0������>n>��>�̶]}��`�<�:�1��<+�t^;}_w��c@4U�bS�GUÊ�W�����ln�|$���უm�}�k�ݿ����n򢭎�iƣ����LhC�3�R]e�b�����=�'���?��!$���͛�$z~FK���^{�%y����֭kr��m���y/ ��Ƽ��X.2fr<��ӳ�����/����D_~�o2�V�.����`�z^/���E]U	��K��+��m�r�	UY��~$US�c$ �F�	CY��m!�h����y�^T��j��ea$V���R�S6�����Z놮D����V���6ŊB)��.RH�"Έ�a��Ęo�����b�ۑ�'������'���B�Z;zX�U�����w���p��M��},���ى͝&�u,�SU�ѫq� j�i�v�VVˢ�Nb*��M�u]�4~e2�+g@�6�L�]' bp�ć��Q�;��|�`g�2/��Uvw�y��w1����,w������u�v���s�}�m��Ϯ�;�\U�{�r�\���5�����e}[Q$ֳm�UH83b1��NF�`�;N�
ׁ�,`N,ʲ<��}�����{�o_�G�1����Ζ�@�7bp�2���FTU�tz��d�]��K�1����*��E��
cW��'"kш5��#��ćh��I�v�-���A}�hR��q��x߅�K��&����Or͞t}�lE������-"�!����bڞ������-t>	�[�3��;�N��s'>�"�����.Z�3�#�{o�.���=�ۿ��F�S�����n<��zIeGLƻ8�}H3S�7�����������3��S�uq�+*�Ұ��.��?�{̷�_|���A��k_�j0fk�����0XW�\IQ���^���*���7ٹ��r�d>�a������w��.���7�b��Ʒ�O_c:m�ؾ�׿Qp��g���}�>����C*�E�
����|�2[[[�E�1p8=��*�޽�|����vY�ZV�zHz"��L@���u]3�1�HF�ѩHD#�}z=���#��xU-*'�d�轧��GBh1&eE���`�*bPE:�m�0���~1�l>}�ҥK����O�H��������ϗ�[�������m1jcۺi6
W��Ъ��^����v����տ3�b�x��A������W����#�o���@ �������ZJU��V�TE-m��Jdo[vؚ�u^���G�~;��33�@G�)�V�h�������j�6�+�_�儉�M�)CJ��z�CE��h�X34"v�Ī�¨1�Ɏ1&��� �1��Hcw��UF�h�NJ)��F�T�7Vŕ��B�
����/��FS1B�9QI��(�b.����c�U��{�1��J�$��9KԈj"��%�?>|��;��f0(k���]1o�{�e�����"��q����UUm�����><��������$�I�[BC�Ӂ>�^��v~mXn�@c�m�aU�@V�x�z�]g�B����|���ĸĺ���>��./�E�r�h4�|��+'4џ�2HȃK�Ԝ�zM�>y�/Z�����BL!#��d�cS��XGaEY��mp�`�T<=�7]	��q&�+�D�U$U�ǈ���U�j�&��Ŋ������CK��}g,���kJ�݂��l
s�Ɣ)fU�U>3���o�"��b�w ��j��ekg�2��$@2��Z��cm�u��^��Oh�oN_������u%��h v,r��p�w���w�������T�
��&4QM��p��S1,+ں�駟fcc�b����|�������m=�G�6�2�Lx��g���a�\�\Ԉ�ˆ����~�����m��Q�>���{�R��_cwg���-�����6�����W��K�N�-'c[�-���9��o�����'��5=�ym��}4�����0�%8���m������?3��W���̋Yc��g
���ǖ�%�,Q�:���Y̗�8t�����n�_�n�AU��h4x� �/^ؖ��-�ҍ��[ΚƔ�T��Q���F5�\�/Ն�YiŗfWd1Y.mٌb#��P|S�2nצ�%���cql�غ��3��`�C#3��c�##�����DA�v �T��0��m����hCB,�ja��0*Dba��P)*ވ��6D�J��3��łE,�(�k�Q��M*Uh�b��(xm1Q�xL4��8)�-�q=�D�U^	�Z�$��hX�c79t��=Fl7����|"Q�JFa2i�ȉ��b:���Xi�t�T��,T�:���Z��ֺ�lCx�����^�ڷW������WL�K��R׷�����~�;�	��ED��{���klZ�N�6ޕ��|�Wn��҄`���?ab<�1����?�hW�ҦbھMu>�*!�T���o����~���;�ۧ@�����3,���>��0�:�x۰�r\7�NV'�Z�? �͠���
����_Ɩ4q�B���U��� �2���d��d4���%�ii��K�6̎���b{k�j8 ����V��ʌ�l�(�#6-!$?���p� kS��������ɴY#8gp��XF)�W����s��G̎8:�&�Zr�zM��ve�>�a�g���ON���>���?�<������Z�=�qw�C�F#��qVY�,x�`��~��s<��|��lmn ��m�x��2�s��}��?����G?��G0��(����cBL&��P_Ӵ5w>�,����W���^bs��h�W�C����#�{Ɠ	M��=>��V�������;n�y@�JWR���ʲ]�`���ɐg��A5|��xBi�Q�BY���W���z��\T�9ӣ#�}�O�ٛʭ[�0ư1w���	�13��9��#(�儹�������G�����l�Lp�b5⌤JJQS�@��h@�*<���(���h�����bkk���.5bE�h2���(�����-�_�H�ث҆�mf�/�Rc��f�����Q5����8�1�oC4Xi%X+�x6��v�q�k[� ��5
�p���'�W#XREK���FBT�i	�k�cpEAT]�1�h�����)�����1���1��dzL>[ɲ(
����MB�iN��(���H�(�����<���x@�%eʧ�4���S���7��z~,�%��9,�n��e|�ò�:a�h��l*-L�Q�vP���I�K��Z�����z�1�V�ê�6�Ν;<��4��W��\�uӨ���=����,��* P���	8	��X
��Т�Q/g �*b�6��T轡��?}�M���ݹĥK0����/�ı>������Y���9�Ұd�q������3}����`��Ƣb��l��8S�6��W�����p��.�I�d8��-A-�i���m�߽�dk��y����y�L��I�;5)�k
Ga,�+hb���X��eQ`]*AU�m��&c2�1� gk����7��$���>g��{o�YYUY�7�E��Q�Ƃ4��@���������E�e =Λa@�0�a��戶�#Q$5����ޫ�����.����q�fV5�ZlJM�Hd޼Kč8���~߅v>���y��[���}R�H���Cj����Ϻ]���ϧ�>k�����c���p�Z�72�u$�X�����֏���c���Wv'$o��C�p��G����-��7����+Wv0�,}��R�m�K�����-G���4-J�O�_�am�)ʂ#]��t��PJ���q/�b	>���������>MQ�� �cL�-����}f�1�g��S�y|� �uG���Jcl��N�|t�.���w���b�]��R�Ӑ��R��/'��X~ު%�Oz�R��,P��5����L���>|�xTR%ZChm�$���,)^|�y��^�g���}k5"
���c��'''j6�G�Ь���!xΦg�m��S4vL�>4"1�I"��Y�8��ql��P���F��Ry�4)��Z&�Y�I	b�q�齂5Z[�Ŝ!�k����b)e8���^�1I��L��
�"Ď�d�QS��&��cDooF���~�1�R����-_C��J��q山*c����,ӧ,)�?/R�$	��N֪�bAb1O����w������|>�(���q��5��L$v�m=�RZ��{��ۇ{׮�ͺ���Փ���*����S��[���~���KӅ�c쒮�Wj�B��4&��Rk����#�e'�%�sw���$�a�i���}���4H�n������h������2[�ns�ib5���>&�|9�S*[�el���i2mC��I�����dl�}��aP�p�7��˽ֱc��_�_~���]�a�V2�J���ڶ5,�sl�c&��{�y~��W����l�R�y���~}pW��5Xm�YJW%�B�ǐ�g��aB���8g|$dQ�����kLF���~�Ǆ�e\!� �V���$���Q�iړ�u_�>��.�o�U�Fಜ�z٠�ؔT�АT��<Ea��-'�;4��t�l����?z��+���r��{��o�?�/�e\e��{��)�fOX!�.�ܑ����]�����]��\�5�_�썶�F%���:3}C���pŘ���[o�g����{� �|�J��y�Z����)�t�����%��]gsm�����h����,jR
4������~��?���Kl�<v�O;.ϯ���mۢ�����rQ�K��sy|�s���{>{��A_�R��g,�9��o��W^��g�ak}�_|���66��>���C����͙˔.��E$,�?�E�0;;e��7S0�L@ �@m۲����%Qʠ�,��Ƹ�{6nY�L) 1� ���t�A��kT0�0T줘mHR�������A�)k@�����rp��2lF;��,�gȃ
B�������(M�l$�\*5��5]�0$��2dKt��yã�]�o�s�=W,�;�FS6O�èIHʙꔲ:I>~ou�7�DT)�W�@"=!�tm��	Nk�LֈX�"��+���>��i$v��cR�h�"�d��y�~
PΟ���Z�f:�L���l�b$�K�D�T2�U�2�s���灐�b3�q�Z���l=�=��ؕEŃy�G��r���X߀Ã'3�(��U�����=8s|Ri�ݡ4�*+�XIL�@m�ȡΟRPy^jX����Ӷ�c�D�(M�\:��a݈�_�%����x��g)�����SG���7�r��u�z����{x��S\f�����Z)S8�����=
ED�mA"���\��~�|�����o�)0v���-^y���%�D�,z�]��	�$$��3l[[[@&E5M��p\�,��� ?����������MI`�j�DD��"���[�u�l������c~�_�����IL*�IM�g\�o�X���e,�AE!rvẋ�}��]q��1ׯ�0����U���m9;;�YM����;��֛|��m���ZML9�D�
�I�tDbJ�2�[�ܻ��ݫ�nl�QtmK0��D
M�/<z�����cP���5-���m�t���@oU�XfE2p`K�ד2}����c�����o8ހwW2em��ս�vm�/�U~���ʋ/=��x�o�I1��r��=�ܻ�b�@k(]%9��B�U��$m�b���6@@���uH�h�~�$�L`L�<��>�ڈ&�{v.E�ҽ��ܨ%��h��!F ��V3�0;�^�NK�z�(aI�QY�{Ũ@kM��sMU�Y��UI�JΦ� *�K;���ͥWb��A`J�y��HKJ$���%��m���zi.��/�����BΚ&�
D�Z��lS�\�>Hv-�]��9��$�m(J�-T0�E��Vִ֕�n��!Z{"U�M?x����x��:��e�ү����Ԡ��͛�����b�C	�AL\H�_��!�����hKf��eP103�Tbvn�j��c:�Ҷ-���d?ĵ���O����k~�7�ĵkW���:�0 �(���%�U��<Y�>ڶ�m�eve�֨4���	�O��}R�OD~^��}f���$��߱�q%/��2�<�[tM�qt�iy��*�:�X���:89��)1�H�cz���`M")A�6e&�]T���c�ꀖ<Y�$�63s��1vFU��`L�}T�5���(]v$899�n*���&�?�V�K��GW]e>�������-��Kr�R;2�~����w�XD����K��`lD�fѴܾ9;����Ӈ<��#���8;��RYJD;K�36�Y����	�*)\)pvz̷��/X[[cT� ��>�)M�55)vLώ89="����x7�=�_�P�Đ��$�ȁT�8�rx|���w(]�����W ��wl���,s���>����$8mxZ�Հo��2(*(����kVE�/��e��tP���X
+E���&�W���˯���̋/����6�-9;;���qp����I���5&eE�,��@d<Z��J�F2.�g�Z��k�L�3�z��#J��l��[�M	�Ǣ��2c�Gi��*^)d̲��#,�g�L>OԋŅ@{(���R"�\�,sŒ�R�ݘ^�h��J�Ϥ���y��R��#�@�ۜY����;��R��,9�Н�\�09x�1,�K��u&� ����H�
LH=�C+��ω,-�͘��H�A���%���)�K�9��DY:�Q�Zg��h*v��	=
^TJ����>|xT��u�vۊF���*�u�֧}}g�!��إ&�i܅�3]�"�EU��}��2�މv9Xr����g���2u]g*�����Ψ�*�y����`cc����S���vy�X�s|R�d�<,�]�-%^Vu�T�da�ՠo��w�?ia�y(�B�陼�īuΪ�!E���v-ڕ����i��,������ѣ.�r�
]�]ؠ�uM�4� <�b��{������*V	��k9����*7�^ac\H4!g1|��NV��*"@� ����~�V�����������}�ٽ/b[�Vk�*9���В��[X<M�,    IDATsF��8�8:9������\����t���+	���f(m�L&�D���Vk�V9!�-��&�LP=�H��ZZ�*JRt��Ih#8F;B�X#9Ќ�A:0d z�$��>�(�)�����k[LPH�>h�{�M�u]c�f\U,���tX������2�N�J�����q��K�����R�i�6��s٦����g�ʾ\��\�C�h4b�^x��ۿ����Z>��>��0����՚�|���!ggg��_�%B�fQ�PJQ�%�;�=�2�s���>�	fYB�{�lV�]&]��(3��țݔ�L6��~c��>�U<k�D2FDHBO��k���s�/%���(T�	1�e����k=D����
�!�#��uuX��\-��1��91$߷�D|.�O���,��]:�Pʀ���S����fx�����x<^�������8 O0���!�{҇��@� an�B�����6ڇq]�ηm1_̪���ַ�_�㣟_�*��~�c��F�I��!�����cӎ��*A�.�S�똢B�`�M$��Bk�B���g��ʸ������.N�q��w1�G��2�89��sݱ������w��z��2��W��g&�	Mӡ�FG��:/�� 채�>�*�y���I���}Q,x�)�H�<�&�e1Bk�'�>0��:|�ΒR�M� ,�g�pq=�M�1�@Ȼ.���b�DT>y���Jڮ��c�J��H��q�1d��s�%�y����/�)���Oh�\�$?�{*�	���3l�bʒ�K4~����OL۠;ێzq��?x�޿���X�1�ٌ�b���,�3��poL� $O)�Γ�q}prF�����f�`R�"����R���0�Цb����^y�����^f<���#f������c�+0�X�P��Ԣ�`��k�$����-	�Ǩ�C�$�ypvL�E�WH��)���s4O�߫Y�լ����l (�X5��Hm�H�s��P:au���)��d ���\���Y��:��u���ɪ y@e����'_�Oi.�����Y@2��.n�FG+/���� ��~�dܿ0�TU@K��[�������5B?R�c�B�R ��M����W�,����{����Q��>���������Q_:,������Xl��q���{��f��L<�nnKt�IEI���Ǚ+-h)ʼ�w]ۗ\=�����lpzz�3�).���L�6���ec�2C>l�677���㥗^�W^a�ǜ||����CX���98Q�tI��ͥJSN0�-�1��Z�����欪*Du����r#�Y.����pơ�b��
EL�D�wC�pe�[��)&u�q��K��&0CP��h��%��r��N[�3'!O�S��F*��O����=ñ�y����uJ	����r$��$GW?ؤI�8�|��1�D���i��}�����ID�d{�e���$��j�\yC@ň��|�R҅V�`��U�k3�ו�pvz�N��֞NO��3ƚ�Y�g�y��=�'-�Jb�����Q�S}7o�L7o�q�ԋ��AI=�L�!	>D)G���$�8;��오 %�C�	H�����䄔�E͇wnspp�h4��8<:�J)��)u[c�S�~�m�����3�<�̦���1��!S��]x�J���jľ�.�a��ߗ變���!ڶe��.'�Ld�����i��6����Bz�=vy�_���b_��[�@�<��rP�:��@��.ι~�]>�{�G|������g>] �6��4�C%A;Ka,I11oj�6(k�AR�@��i&��gM���&v�7���T��d�aM�i��zA�,�E��(2�ue������Zj��&���������o���D�2c�$��z����R�$�p��h�$��gQQ��(ML�#���XC1Ҙh3x\G��^J!KH��AZd�hⱅaTd1���������)un�vy~��۶���ev�m����M���Ӵ�VU���ll��t:�����9��������UU1���2�N���9�������9���@Y�,[N���H/�;��$�C+�1M�\�T�5���!B*M�µQ*c�SPK��2�ѯm������,^9Ɠ�<{Ѵ` Y�b I��H���W��(�Z-�'�$b8ߘj�2�^�4EAY��ev�ϡ�+X�,�f��H�xR���������D�QHt�H�.�XIT�c��pI"�:�$&�5�P.��M������"�����J�$ҹ��l{29�R�#J�[��O�yL]gT��k/�S����w��(�V|S��1�&��t�]B��ipe)1&e�5�+2�8�Z�v���$@
W *���I֧�֖ʍ�WUf���(��o�������}�Y������1fyc����KA�%-�U��0ПTz~��-�N���?��؞Y�rY.w�s��A�H.�̯�S��L������3��"�i��\��dw�����9>�������T� a������os|4�t�;�����A�+U�Y�͢fT�\3�k2+�B��tG�����A��L�ߚ� )0��Ѩd2{Weצ}���C�/K�1��.w��)�jV��ṡ=}�XeI�u9�c�J�.�B�&I��8kp���U~l,�p�a��jC<�u�"^Z�}X�v>g���j��	j��E�l���A,ZU1��Ç�<�LC��UÆ��nX�{X�>�~���i�~��KU�O
���Cw</m /�_��|��5�ס|<ظu]���׷7��Tw�&W����&M�pxr�$R����3��E��mhЩn�&H@�E�yO*�ULA^�R8OzĔ(�k��Q)bL(ՓP�!��+Eˊ�P����}�ߺ��A�֚�u9�3�a��ƈR�IU]���ka^g����>j֞a��r=��X[,��(���\��g��\�UP���(P:o���m�d$%�E`:�+�-F㔱>�wI"��PS��Ux���N��Y�1Z�L�ԑ��Q�BJ���4����8c�c���AQUGhӖV����%^�w�o׋B��>�%��hL|ԺU��wQ��s������w�?zp��Ͽʯ��o1�w�fZ�I%Q"����.0.
�Γ��gKfuM)��x�h4BiǼi�ǜ�f��_���)W�^�C�tX�2�vri������3}���Cv�I��1���l��/(�vZ�#(�9��~�kb̯�:I��)u]/�1�=���ǘf�%����K�x��jИ��^��������&��[���g-��Z���K�so��]We�����9��BYE�	c���	�g� �b�T����U�� ���F��>upp�|:є�q��с�DY[ۦ���Jn�f۽m���U��O�\���KV�gi&���� ��v66؜\gws����̆���}Y�˟aR_��2*�Dl��i�(�
�
RR�ń���L�
5Ei�!��g�[�vX]������{�?⭷�����dz{�4d��11��$,�?��w���\�/��Ļ�T�6�K՜���0����d�����bY^�_��<�y�2��:㇇
� ���0�/�����z��l�9����|~ڟgp�4I:�Wh�PJch��}3� _�����:��F�eY�)8�L笣g�d��2�A�F����g��� )S$a��$�r�f�-�%8Pl��QYĺig�^҅�PBt��b����F��8|����eц�ۈh��s	9j��eU5��<r�RI�F"��)��ژ�� $k�Kb�(ZDy�@C��AsY��A:��� !�4e�C�uRZ5��F?&Q *����t�Gڮ��,�WZO��b�>��?9>Y�����uk2�|tvv�nݺ��������o|#Z�tA�mT��:ejچv��Ç|�{�t��ʫ_E����5zM¡mB�'��l~F�8g�eMΜ ���{��Xf���&J)n߾͇~����:��e�(1�zͥ 	gt�>擤/��S����o���v�)KCJ��K�=�G�L�ǘ�a�{"�Tp�s�]�y�
/��I��j[�S��˙B�;��h���N���1>Y���T����J	Lv�2���+3OR�j�h4b>]d����&�H[wh���V�R��O��:66��~�W�\��m�J�A�Z�lIQ�K��#?��yd�(����]�|:#t�|�����*D�Y ��(�}>�W�y�2T�o���W��	:o������.���U~��x��u�no���Q�rR_��iU�a�,��/7��F(m���^�'�6�����A��e�ch���܋/PM*O�xx�0c1����z�]�k�r��t��_���փ�k�Xt��@�B�y����[Y��*���`p�?�[x��o����:�Z��1�u��Ou��lvJ�4KG��k������nBX�Ƙ�n��huf5��:�?SBʏ��X�eV|r�tV/��j�`�!f۽\I�Rk"BL:����%9��1\3Q8+h��&��ߡ$W(4]3mU	Y1YD+���0�(�E��*�yH!%���䌨:�&���耊1�d�$��1��Je�B�Ť6�W���c�7�R�Q�R?�H��� ")v1�n4��z�4I$ň�DItZ���Q�F���gWRRJ�N9R�)�@�:��EQ�RJ�`��6`���F1���c!Y���=|l�����R,�v][We�������#�M��������NO�)���͛	mۦ(ʏM<⵱�j���x||h�|�Mv��g����]��DaQ�����ʢ�����|��tF�����(f����e�w�L�X,|����w�_���q!K�m��檧��Rͽ��0{x4-���'v=��cT?��ˌ������w�mH�L���������K\��1/�D��'�<�W�.�Q.g
����Z^�y{��Y��N_q���1�Q=z���&k#�ɓmU�h����d'�p�j4bwg���M���I1b�e{k�kׯsew7{��`|��{i�~F���ǿ�5=z�3�6�еs�����C�y�������>�ڞߣ%�xe�	)���|�?��b� ���3}	MJ�-*����+_�*���*���6��u7$\,���q��φ�M1�2�"�{HP7�B�P~��ӏ���@��w�;Ϛ���=�}�y��w���RYn�e�>��>�|?G0��U��g��n.��9��Ԭ�hV�g�˺��dyNC�ou޽,[�j��Im�����ܝ5/݅���������_���)C}:NNN�������l�����X�0Z���Y���|���6%"!%��m��`��$%ڈ��5L2F%AG笏	�V��*{�)QP-� ���Et�f�����[��$*DD�GR��9E�,E�����:�R-�)Af�譈?NAG�t��L
!:e;�z�/Ԧ��h�{�:01F�I@2�e�Jr��Z�C,�1��ڤ�s1�co�E
��>����AW�R�q�I:oA�l�K2��Ҵ�b1��8U��Fb�֒��|�:b8DB�	�ċ�6�I*��T$�BE��`SLN}*��[��	":F��Rڥ�x\� �t��!��HL2���M�
��Sw�y������w��6��|��.����.�m��|h�G&���j��*�M��|t�6��o�M�s/|���7pE��]h�� ��X���1�o���Gw	ƕ�MM�;�r��ƣ��w��?������׹u�V�yBJ�΢�.�!�C���K$g&��T��x��d��^\�.���Up�jau��9�d0�l.w�������W'�U��LG���]�Ւ>N�>wFY�N�>S���/�X���rPk2Á�#m]s���x�}�]�P=�E�ޕ�dbFR0*J6��xv��n쳳�E<"���2��I/oQ��^��!@%�U\�v���u
��8���7x����[ob]����V���=���f4������c��Q�K�~��xOkB���#�׷��ڥ(3S�	-�"����Ĥ�*���9�yՒqh�Pt�'&ͨ1M��UD��ʡ�%r����MP��Y��)K����mP��t$��-�t�� �3<����'a�T�!����WH�l�;��Zz����������w��t�z�u�����r�
���<��KH�q�����ѣGܿ���q�-���$�]�-�"aHQ0�����^}6h!6�	��]�6�4���?-���v�)tSRH�ke��Ց4Ac�$ʞ�������"�nH�KI�Z�H����`;���`;��N����L�T�E<�v�B�Z��C����͛7;��7o����������YF3�R�r�L�Ke��t�m�Z���}-B�)�I��6Q�eT2R*�]J�������_��$c��H4��N��N�C��%%��(����T���1XM, M2�A)���D�26D	$/1��$m�^Bx��,=�����VX�'�R�(U)cJ��	�^D��C�����(�]�`'6�-@��zܾ��k�֭[�d2�����3}G����6v�S��o$ԕ�	�4m[�빤������������7��ۿ�;���L��P"XWr��>���ͭ[���{[R6���zu����$�s|�]�r���-r�>��7}��;�Y�~�����|C�u�f3���@�x�JXH��f��]N(�I��30}VŘ��1����񒲿X,��j��
�]=��.����0�(Q�}1�r��c�Zf����s�RFH(��җ0�����6�@�iY�0��[��g��W��E��#���l�<VVWJ-˙Z.�U����^�!0�1�
$v�l��W�L5��|����>�U�{'���ccc���X�M�_.�>1���-3n}C���w��7�蒔�.%*m)ʒ��9M�,eo��ˀ�+�,)1�ϗ:��"c�����ym�����F�|^x>f6�q:=#�fm}���/pew��x��rL�\JʘMG�.�*c�zŇ���/���6Ta�F�
�x���Pn,ن�v �V\>k%d��֋Ռ_J��O�I/��h���s���>�^�h�y�l~��"�*
Wa�Ba(&%����`}�J}�O���ƍ�!&�x��G��sաq������x�"g)t-:"�4��3��d�>�L i�L
t
AGҺ�`Bd+A����I	�(I��1�h|��jQ>h���n��u1.?H]���k�(#���o�{���{?=��o�M;��IXخ1�ģ��Ye۶momS��OZ�N�k����h�8��W�0A�^��A���(���l�>�N���D�2�����$��BҺ��!im,ؔ�7J�����	ګ:�dt��+���""��:"��d�j�H�jD�����dc=��1�%�-7���a����0����<�G��>����۶���h#���;j6�����GGGR������|����g�͛7���3}��ݓ��BPb��]l�J����b���,f���G�l~Ʒ����s�/��2/��_��Wi������_~������t�h��u%m�b$��'�����#&�k4u�n?��_������]<x���d�`:�����l6G�Q5���O��Z>0=U<��[,�e�b�^<	�
�&bub(˒�|����d�s���A�o8�����R�X��놅�9G�$٢��	i����%��i�[c�f�R�=(��m�msV�y�-��tߧ�WK�O��i��ӊ�|�5��|�<�sד�k�
��8g�b�ʒ���Zm��l�0�,�:fӆ{\�,���(HQ�7-՚�Yٽ~b�(
�
�vL��''��*~����u&�1g�9��#�lsT7�u5���=��v�$�,	m̦�*�G�N���V��C����e;D��"!$f���`s{��G��;x�w�}���m�4UU�������b����a!lb��Y�k�5���3{:y��9=;�l6���
�_���wx��W����_Ѕ����[lo��}�m<�zE�hpnDJR@T��������S����.�~��=F����2v�r��c�\��kw�A�]n��q�u�1��ʰQY,�ι�Fί��z�j����������3�O(�x����׾�˯�o�q�۷?���^0����sm��    IDAT��Õ5�*{�lf������Y���U���xD�^�a4YG%�(�����t*v�(U8�.�+��קg���zWD�[ԋ��h�����uR��E�I	-J�I��:�3��%CM��E"mЁS�T��̕R��:��i�ME����	�ES�H�֝E[�u�Q:c��C�����d�>�w��ƍ��t ���tW�Wڣ��SE�(ڮR�.��Sl�N��F�I��騬�$�7:��ѕe�&���]���@Yy��EQ(����Z�ԳL&�|�?����1��R:�=R���c[��h�(^=�1e[����.�2�m�˿.���՗�y-�z���y�f��?��{��{I)�I��^�"���o��7oݼyS_�~]'�nݒ��뢔:�_�D��g
�nܸ!'''҅YD���6F-�Hl}}ipP�Řӳc~��-=zȽ�w��	���r<��v	�C����� ������g8UKf`�u��o�{�23��/C��U����Ռӻ�1 ᓹ0����m�Ռ�j���`�z;�2�0��`��kX����g���y��rPt�=��)�l�_f�rИ����8������m-:���rlݓXW�9��FL&Fe�f�_�LҮR�eT���Ễ�Z����Y�(���p#p���!��5�D�Q^~�+���qmo'��R��jD�\^�,����Υ���*����瓼J}ILe�Ӱ�J�
�\A�f3�Óc�z�-�����0�N�ЃA����,��Z�2�K�
?ϙS�h���"u3�mj�7�4�C�tݜ�4G'3NN�\����~YS����[;lnoѶ_�%���i2�{P��E��T&(��ڹ�PyY-��*\�/�jyx��q��Bsf�Y�c�7�{{{���s��RJ����0���e��5�}�Y67�������N3=�sp���GG�����M�)���r��m:�2��u�s)�(�N�ֺA̩��$/]D�7m7&�p>��a�����]���C�d:%�XGm�B֊�l������(������H��;���1&km�˔�6fjִf2��Η� �@g��Y�gG7n�P����������ɭ�o��o~]�c��y-���O����h����qP����p�{o�븷�'��$����w��ٸ���' �׮��\����]������g��6����n"J)�7�P���������͛7?���)�X,���RlD'%)���(���$�o�D��}ĝ���޻o�������8�k��Qe�ۚE�bBi���v.?Q&g���
���{w�����RD[CL1냹jI�0.{��<!�A��qy�_� ��eЗ�;�hm�'�:R�e9�^�����~�iJ	���P����.g!WI*���I�ße[e���U �OlI=����+�(H0��'y���Y/��'��y���]}���V_Z�,�٢��8WR�2k�T�ƣ5l��7��D1�1QY��l]�!�^�[����9>��Y	���H)��_��:��rA�S�.����1]����J���~�o��ݻ?�������V�uF�k�;�`�B�\��|����<�Α��iO1�a�1(�����^f:��d��o0�����C9�I�h���E��mO�k��0�\� �ɛ)�Կ,�b��[�E]%nmu��Z�}��.��������[UU���q��5ڶ�?�w>� c�Q�+ƌ�&��g�n��3���w�srv���U���_���g���Z2���G���T�k��{�#��]�1��^z1��W>%E���
>mt!mn͛��jT�%��֣���6<x�+��N�y��jp�IT�Ϸ�op��?�� �������F׫�t}U�8;;���}�5d�>Y �)��g?�����7�xC2�J$��Q֤�bL�ֽ�M���1*K�QI�����p����[뛘�Q�����9;�*�0��l��*�NO	OY�Q�}̥7��!P���|��P�a���<z4������� J�����뙩)Y�W�=&*e�-ԋ����A�!?o��-�x�ؗ���x�s!C�	�P${2�~`�e�J�(҅�����h���^ �|�sQJaz�R*gy���������-Ύ�LOg�U_��nllQU!>��$^�#���\��*C&���4+��
1�",�b<-�i���RZ`:mx��i[��<IV�|���2�'rn��9��z�ؕ�>E
��(ʲ�p���<zt�ՀQ��DSX��sy��(����O�*RRH(�}�3P�&��FkGaRL�$c�E:i�@Y8��z�O�l.K��-�ۜ��E�{����AJ��b���1[��e\Ul�:�O�sl�@��d}ס5M�o|,���lll���ѣG|����3d:������!�����uR�|�+����a1Ei���C����޻��7�}���3f�:ox1�6�c�(KYU��UaݾR$��6!��� q3i�̨��iqf�']�����a��n�͛���-�߻�JYU� ���w����g��q|LpN��"u&�h�
� �����h*�-ZB0β��F�����@�+�J��q.��*�J)NN�X+6pz��-�T'''(�;v�#m�E���O����2鳢Ö%zE��w���%� ���)��y����TB���%&��5A]��w��%>�]��]~n�g�L&�e�R��%i���l/L`O._|���P���"*�%Ԝ��F�<HްVe�h4¹\�H�H�@MR`KK5���� 
��r�o��\�g<8;ʾ�"�q���5�5-Bbzr�b!�Mã���[o����%������tn쾴��S.g�SʎO"�|^m��}��^�AeW�k|hP��h�$!� ��e�TE���d}}�Q�G<XMu]G#]�)��͜z��ʻ�esͱh:��
0��Jh�Qo]��nyl�5�:��>����E�{�d��?����8;;���l�m09����{�fY��L�Y.3�m{,<")I�I���g�{f�4?�����1׼��ŌbbB���H-��I��-�f��X�UY�l�� "���Q��ff-��{�w�I]׉&�U����7y]����#�ׯ�tp�.���>�p����c}��tzH��3�N\�e���C�ܹ����{�pzzLU5vGتi��`�A�H���hă�cbJ�G�x^!�Q��NC��EuX����Q���?�<
�|j@��NB�a}t���ѻ}����|�HS�	O�ƤU<1ZF3�/Q�����R���x<N�u�\I ;m��9��Ϭ�两�\������,����O���R�g�.Fp�c)�/ט>����jR)�(O�վ�h����%ދ%g�� �]خt���:o]�i�T&�d�£���v�.����'�ː����^`�Y�]Ӭ��Nd�MSqr�`Mz:f���;�(
��1{{{���S�z�xx\S5�`��+��ٙ�a��,K�����O��_��=�Ō�}���)���%BF��P��o�nS���$t�o�\)E����8�`]IU� F��A,Fl�vM����ʵ��'�le2�"g4����d42�QB���89z���}�R�p:]a�!4���\K����I�_�1���2�ߺX��?�?��:�,ĨX.�<x��g�]gT\[$w��2�֮!0�5��)[.���ײ�i�֐��4~-�������,������l���	�gS�k�Z(��kCʸ��2]�MK��v5&�8�PRJ��PR*/|�Jeh\���'d9�9͏�<���N���!�\2��9+���-uJ�k�����yCp.�]��191��X�d�\�Z;�L��%��9�Ʉ�d�JFy� ��j��I�n�8��5z��)K���6 ��������^b\��&��D�&Zǣ��me�mj��-�|li�2�I������j�|�Iܔ�~�Y����}��q&#D�!��uBЈ)˒���Ez�
()	�1_M1�0�p��^�����:�@�gU/899����_���H����P�9�k�9Ҍ�ӓc�}�!}�!W���h"����2��dNc�o���~��~E�����g.�\��nb��`��x_�l��p6)�Ȩ�J�ɜ����	�W�GH�qu��!j�`<Bg�|o��d���=2c��s�w�p���rNc+�/h�ckAA1!�;�kZ
�wTU���@���[�D�x��:~� <���a'y���$��Ln֊���u�8:�������J�RJV����L�S�s\�zm������'(m8=�rt|B�8�T\��E�L�g��2�� �Hcc�Z��I�=�Y�j���*�R"e!6RHʀ+�@�΅:��%��zj�Ş��;::{{{ ���T	�*��2� B�	`�~�i�7�c8̑��r5c6=C�W�itk-�'5
�R�}U6���a����畗^�,K�?}p{-q��i�t�۬�I�M�ԙ�ni�;s/:}��]��8����1]V��j�M:�"2*NϷ������$��R
緛5:G����OB�O�������N�O�=���c ����ϑD�b>�SU�)��i�b���LF���|�;o��oP�%���ܽ{����/eN�S����#v&;g�������G(�2����lN�in\����1�q�n������'6�9�_:���L�����8�D�J� �)ڌ�a���8� Z(23`r�͛7�Z3�B0�s�sh�s�{��x��!�������x0����hA�I�$!Hf=߈��Ĺ��ŝ��S��~�ƹN~l#���]]� a~7JJ}�Skm
$~��}~]���hKʉb00�毢(BqrrB�0f�d�f�u#���!�̉A`��65B2��,M���R���qȤ���h!�*�#evp�ɫ�<���yjP��ʻeB;'c��e,Px6Da��%�w�P��L�}�&ZJ�U�'�%:�R�I<���Q�3�_2���]�>�`4住�嬪�=|-��6)cb]D�ClB�'��rI=O�����
���T����đ����k�pEA��5�sG��F�v$��ш���ш�j{>�Q��Ӻ�h�}� T��ު�X*�x����g,�(4Ҥc�
z]�k���ڲ��l��?�l�IEuQ!Q�(-p? 8�My8;c�sA=A@f4�ȢT�N����⫯����{&�n�w��#n���g:;ag8�����OFL�ƃ\K�.�$�!2���|z��l���c�,c|x�Ji�޹˭[���ڿƠ	T�$zEt��j�z����mÑ��T����!��L�a!*�9D��	/(�%�@
lA\�`�O,��rF��x�9?�1�FL&4�������r� %���&3C���hF<c�L‸X1/�I���,�r�w�s>K�hw���H2r)p�$���# �V��H,�� �D�$b@����}ָ�3�!S��@��Q;Bw��5���0���|�n{�!���$�bIPK�h�*�W�*g�<#�y1g:}H�^چ|�SN�����BtT���e�(��b�S[O�
e
�R�& �%�Q!��3Bt�:˩}���=_��tӃ�(���dY����D$���HU6��n�7&j!ڦ��$8�ɵ�6KBY1���<�ލ��[����-�Yt6 �o��&�I����q�h������ ���"�k����f3vw��9��)�$(R@���]`��3�ZQ�"8�$Ǧ�J�DV�Sޛ�L&��^F�U������ů�����6j<��퉝>S��j�@	UAH��&��QV8��*z�7 �l�	y!"o��C���minUUF#ƣ=�v��ptt��cM/��nӤj���\&� �H��������~��G����˲�����k;��.��W1������$v�4������Ͼ����7r|�z!������CU�h�g��Wi�o����ۿ`>�!�g0�����,�GX.��eI�u����h{��t<��5�����y���W�\9`�J?�֯�K�])������֦_L�9Q��4�"]M��ԡahr�a��8W�G�4�lg�f��{���U�9���W%���e�bV/@�)vwǘ�yd�ne��@������< ��Z��)��5���p.zdLk�T�kc�U��/�kO�5y.@i��8"F$�t�<�2jv�;�U��p���b"�il�ZЙA��R�Ň���<O��>&̥1
$R�q"uR��ֳjV4!$�J-1m�'Ĉ�ms\�ԫ�S�YZ/BXBk�R���;�p1��λ���y�|�XϷ���l'�"��2\�e�/V}��ٛ�s�9��9���l��Fu{G����kmn)H�TQI�P4v���{��2��T*SR���u=�|�X��ƞ��{���ѻ�
#Dp��"�=+df�RB����E1�v��G�m�VӀ�bU���!5e�%�.K6�N9=�1�9`<9��uP�����-�K��[N?h1֦ITV˶SJ�G�G'R���1�;�q�Y�&h"���7h�Q���d��o�
ߑ(7M���ҿ~����E�b+wU��e �/��ߙ�����r	@����C��������c��1�6Y��9?}@9��*��\[/��s��"u�M����s�!0���4qgH 2�s�R͖�'D���;�sX?����孺��;��!���!�#���_� U@�
�'R��Uę��<n$�c�ݣ#~��[��V�ـ��T�"g.T��̝qڜ����n����oeZK"�y��-HŰ0H�	Uē:���⃇�2�)��C�����*b���$%�%F*D`A8I��Z�:^U!p���T��(0*���A��o-R�����c�Xy�SW{�]&�<��B"L�.Fh��<;OA/��L4(�Ur�$'ELNgHN>���1�!��svww���[+]����0�۶%�W��3���4'�1���>��#�=���N�&q^J�W�\a>�o�/Z�p�{�/�n���: ��ɘ�k!�1D���պ�
̞`�>�/�=Y���M���>�D�;D����2u�n�)SYJ�&L7n����:�"DWR������J.g�3�=<b��u����Өk׸����f���n�2��D*R���.�B\�~m�bv�q�C"�l�1�7�C��2Y�l��Ď3*�G:GNF�e��+�/2���:c}��kj1Fc� F���>��s��l�[)�@lȆH]-)�!�������=�����L�����{Ì�ܠ��0��鮵�婔!"�\s�3"��ݻ�99:�D�o<��ݖ�$�V]�b�h��k��󰋍6�c�����XD�P9�,�RhS�3�E�+3z�`0�Xc��ݵ|��?e�w�����7<<=&�$��S�{9���fF�*qN2f�������4n;\�w�,Ө,G��sM���yQ���GȈ1)�Y�{�Uĕ�L*���E�"ϱNPVZ�LF�lE]O1�K�RI�\L�EA`����
�R8�q.2�r������n�geK\��ZVh�8�z����gܼz����h�T�� ��#�B��1zD���3�߿���C�޽�r�Ļ�]����k���w�L�h�c4�`�?���>����E"��ߵ��گ�\����;���;==�z���A����
��ړ:��F���� |BHC@��b�O9|�ڗԞ��;�ʙp��Ѝ��P"8?�2�w>F�4V�V˖\�я�pg��S�?@*[ "!RElH���p�������egw��xD8:��kB' :�#�Τ���z���э�bf�_n��>�OLj�2e:޸@rchg^��2��B7�;������4Z��t^��\!e���n��2��{�H��Oc����6*+��	�Z�-8���9<<\ӽ�"�h!�D"AK�̥E�ͺ���+MUr�{����!?�J���{RiI��*k����R��������(�!�UJ!�GI�w���`2��4(��%"8p�ipq��5Ŏ 7�|�
_�����GGxp���3]���?����P�cM�H��=�    IDAT���n�xE�Tq�o���ɇ�̻�-�Œ�p̍Wy饗�FL&��4W�V�")Y����C~��=��KY@�^�C �A#<s�Y���H5���6����bIm�i͔R��L��2a���|��_z�o|�ufƭ�>��_���B�(W������[���;��<����
�Uհ�b�m]�3��Ղ���srr�·=����C����5��m!�5�2�w0���N�[�_�H��wN�Ex��&\�)�J��ck,nd>����I�N��.�~�����w|!v�����	t�&:tBB�T�A�����}j{bL��	�BB�2	SB�]#��!Ɣzvn��]��!�=e'�.Z��$�R�0��Y��g=<e��&�`��h̕+W�}�>ժ���,Z�.�D��k�U:�ۍ��e��Ob]���m�#l�`�d�Z����u����T�.�-��w�w?��]�:%�v������וտ��9��Z�X/��k�s�fZ����~5u�VU�b���Wc14H��_t���!il�Ķ�Je%dj`�W�~�:M���w�t:%��r�D�D��[R�.�'�6I��TyW���D@(�(�D��A�;��˯��3�p��!7���rq� W��8?=����4u��+�1�����������sL���e��Q���[�r�`�Y�)_���>�xƭ�������M�1�eXBT!q>�\U�u�x<��7�ÿz����⋘�%ϳ͜��� ����|�o�zĭwn��G�����`4d�J�@��������J/8:����ý{�x��!�yb[�PR&�h�B�и �������o�g��n�,���)�����#������_{�[��_A�@��� �4HA��פ��5:ӌT��9�{W0ِ��-Q
N>�ڲmj��`	�!Q\TU�^_�u�v�����ԕ�ښo}�oB�]��l=�W�9�R�u����-�-��sP�ր֤L�חL�U@MgS���2�H��1z���O1t�ڗ؞��[,�x�J�[�d�B���E7�ʄ��.�'b��%��s0���	���$i�Ve����墂��b4���g��}��%�ѐHj��Z���i#X�kZMδ�zo[I��2��i��Mꮬ�N������m�GR���jM �9|��u?myW���c���x���,��z���1�����S��;�Lf���z���1Bi�ƒy����P��%X�6��hLQ(!	�b���Eƈ��$(J��:�s�������k�ٌ��QK����r����߈����Fӧ��z�I�� ���_��^c�`���r5%�$":�w��SN�ψ.�O�|��-��w8<�x������7i���${�=�����0��x���woS�#E�ɖ�����<��g1e�����7���7��������?�:�u2"�@L�m!�i�L6��3Wy��7y��78ؿ��ܾ�6 *R6�*�����+<��WPz���Y��o�M���3�F��V
��6D!�A u�x�
Wo�ȵg_�@����F#��(oȲ���.��(r_���HzM����AʰY穛����:��/�3�"x�ώ�!bׄ���s�O��W�Xc��*��u��sY�o��]pĺ�#�D�}~w���n��7:���,�(����6@�؎A@(ك�D�w"����E�#j|X���a���G�S�C�'��9��P!(1�{�BJ����#{��׷6��ðvH:G��,"H�ሽ�k#\ erbh(˄1��6��nk�\v���LW��ȑ�#�-5u�nFD��EI��庝e���e�ēX�p�6jO���ڈsv��KY�����A8}�sk�{��*�n�O1�I�g8פF�Lᚤk}��+B ����x�͂I��A`2��/8�M�5�
��(�:�mf����HH:�&�_��8�5f6l��TЄvSsM$7��!���䭂�PJs��*�kN�Θ�N�Ww�yx�Ã�P�h����jQ��FF�_�kO#�EI��:{�Ƀ/��c��9�����������?��]��������8�B��H�(����X�\A��������A���w?��)v)kO�z8$O�"wv��wߢiQUMҝ���f�NNg
Q���� /2��9Z)�,#xP�h8�ȇX/�JB�$U.�w<�l1�G�lW ��mCŀA> x�=8�瞧\Έ��*�*P6�c���e�J%]�G��5���y�����.VQ��6�0m�O�܇�tkS��^�\(����1Ɣi������3�jB�!��R3��-R̤���<���?�?��O���+�R���e���4������j�r�RZ'-�NU�&�~��&V@ˎ=U�\���v�%A$��PIZ�5�����&+��; �8���2M��ʵN�G��n5{/k��;�}��s��Ɋ�H����}j"I�ä�a�j��!��/�[���b�.Cv1&N�~)�"�;�����6e\�"����Ν;��x��g���4���3�s���>�T.�]�wL����>���������>$)ѕN<B��nQ$�b������Ae)�!Yw�^�ʲ��:3�ImBH��&�� ��wB Ed^V�,'8:;�t6�iB$���b��p���$�k�Z��{O��Ɣ����-o}VB�;ɻ��I�`�eX<&����ٔ�����6��}Ϋ�(�d����>É9 3a�г{�%n޼��sh��46�E�x��`1���ѝ{���_��1]���`=VW�y��}�`�[/+��z~������-��9�7<����o�����v
$�dgr����)�,/�^0_�P&������cr��U�`r������hYq6]@��@�Vx-��N�.Ғ�w��y>����旿�%y������b�Kդl���.�:���k7��9�iq�����x�`�Z2��������֞w���_�;���]VuEVYFӤ�%�b<�p��Unܸ�����կ���Ͻ�p�qxe�����V3�R8�BT.dĻ�;��:5~�!]�֮)�֙�6��>im�@�{ t�C���u��.��e�������>Qs�9�:\��{C?�fah��HL�*�t,]0�g�iD�"6um
�����j�T0��� O��?{"��j]�s9Ep>z��QH��A����8��(�E�ڢh�l�ƝgKf�����}�$ӻL&�����,�+�!�QjHJ�z۪2�-�s�Zo��.ӷ���8]SDb��Қ̨��iA�En1b��`P�)q�rBQ�F��d���j�X�i_҆u��7�R&���p�^��uv/e(?^r��e}m���؏����?����M��M]˛n�� ���qHi���̴�w*�����[7�w#D�m`�/u�$���rU����w��9�fMC����v�I)%Zl�Mg���i��������CJI�$AIVJb��2���i�����F`C�ɑ\�Nvp%ӳ�Um��$b�sD�L����Ղ(���,�*GsAm��d�g��R����?{�-��ʟ��C����O�ۿ�[>8���4IUF	B��w�ի׹�ʳ���<{�r1D�{�7�{��^x��_���&F�C��@��!#�)��y�y�կs���64��,8��dʉ�(����'/,1��u(��)��[������W����LN������D;2�Ny���w��ZK����x�eȇ#�!"����g'�������q{m�,ؿ��}E����Y��,�J
��w]�����C$:����������b n�5�������i��-���C�R�*�-�K����#�'o�^�h*�(D\;-���!D���@�x9��B����_�1�D$�@���℻YN���s|������������x�x��;M]R�UXwe���EX�Iڟ��c]��=ן�J)��J
�4dENn2|41R55��$J H����qC�9}��uqx�����9��x�~�:�Ɉ,�Ę�SG�/m\� �>��!��E�>ٹwc��ߕ����9��f��
��0�nC�%�<C�5���q�u�y��y����"����J����j[�^g�c��GR�����Š���\F��T���L�04,WV����5���3�v���!r�`MRJ������Tu@G�S(C��b`~��;��z��.y� �5|>�˧����\�k��&�n<��|ͽ{�����G�߿�(˚�jh|R�@hL> ��q����u���%7���}��p���ܸ�?{� ���{���)�]�j��g^���9w���W���4h-[8�!D��Q&.��(��Ӗ?/�_^V����_��=|�6�|�@��B�3CD��<�V��lJD'꫱���L��A��~�<��V��.�-�'��n�e�,x��]t�.�/��J�����k������[��o�ɤDH%���k��я~�T��Ȟ�髚+"��EAĐ��ZA
�]Kbk�[��µD���'k!"	�sOF���h��s�j�o�x�����s��Y,KWS�U�4U"�\��&�`��,C)�`4m��M�[4�z�i�n$}�ņ�9l]3�(�K�LF#�Z,�d4�v�ȱ�>6M�&�����E�q���9����}�\��0� �+������r�.R�\�*u�_��u���c}'���k+w���%�&�� S��V���µgO\g
A���L��A���(|�px_�뚥�(�ϧ��۬�vA`g����}(A�w�g��甍�llt��Ѐ4�)(��;=!,O8��M�h�9���wyNe�H���+�-.�Qx�8Z�yx^��Ś,����p����C��`�f�l��L��QJ�1%	���J~����7��_3;?&�
�cq�������d~6���y����׾J�<����89:N�6F|��4D�� ���T�^|�?���y��w��f8QV�$�%E9-�xޖ��ylD�{D��Q��*lY��d4��j���$H�9R�hr��8�s�΂I�S��9������H��ҙ����i������]�8v��u�����u��e𕋙�K_�A�bh)�D� �U��Z
IPR
���R*ɤЯya��˿��ŏ��/7U�S���)2}AHQ�c�QDA�!D�Iʑkl���^k�u�.()pw�12E5K���)����W���=�����n�\`/EaA`L�p(�~�()l:e/frB�(�����s(18��&�w!A&�#%"�V��i��(@K��
-����[,TU�sn-�V׏�jO�uYî��{鵍��Ŏ��ǡ����vI�r����u��~8��l��A�ׄdj�%�Y�]I�����I�Q��J�nJ��9���!�+V��Ya�%מ���4͚���%�si@�yY?{��w��(|ʸD��5e�����^�
����3:[�%�����ūe
\+�pT�(}��5�l�K4�[�0�K�ǣ��h7�S&��^�M6��	��g��������;w�cw�">�4M���Q�&7�����;_Q���������q<����z#Ā

�2DTT�����,=�p��n0��?��?}����6�H#��k�TD�Jj1�ֱ􉛲�4��M]!�G�$/3F��B������f�'b�� IXJMҠ��B>���|k�ɞcwO�џ<Hl;�k-��!`]�K���8:�ʶ�ww��n�����\Ƙ�|b���wY�.����(��h�
�C����S��̞h�ԶNٽ�VQ pi�ƶ'���=w�9^��:\����������[bg)�"��>~x��x�`�q��3�	��ٛש��:[2�mCpĹM'U�	�w��~�i�JY�N��{]7QzD��:ӧ�a4`�%�e4��,	��(������lFh9�V�!F�њ�>���:���bЋ�z@�$�-��n�J�� ���i}��Q�sS����uI><Ew�!D��0��q5Fzr�6�P/��S��/"MU�Ɗ�1�>��V����od-^ꕧZ.��\�ju��ޢ��6�,�kb�����TW�o,%O�e���d����>68۰�M�e�29>"d�!�Т9<G�S��y�:�gXh�sc4�h7Y��������]>��`A��DR5�5��p��-�L �%Kp��^$�d���AX0;u����
�
��b��IE�"������� ͐ݽ]�S��3&;{|������]�y��N%T��T
h$G&'�L�J�J	�J�F�Nv\�W-�MIaB8P�Lf������9�k���C�ȇ,�%��]�Ԟǁ��NT�v��>V����`�7Y��z��3��ه]t�c�;�n]�	��˪�� �����-���)cZ먢���XU�(%kQ6'O:n�ڗ۞8� ��1FA$��)7'.����.?�%Ȕ�=�{�=Q�I�	1�K��6C(����ŭ�����7��7��1���ӣ����`�)Z���
����t�����u�|� ppp��k�о��r�!�ј���6�u�b6Gg�"��;�gw��Yܻ���(�+>:�s��ݵ�v��ԕ�����l�'�.K�}�sc����MRlH@?/뎫���/�eY~,��]VnY�V�.���w�^bDӠ�F��5��d@�2�����`?�1�����Y�is�H&�d³
5"�(,Z��=�b�=���qk�ZC�L����������ن�G�޲'��{�#±ZN�)��J&٘���E	�Ai�򎲶(Q0P���t��Zy���<{�G�;?y�����ǈ��/:�oU-��U���܀�+f�#�� �BD� n��,�MI�a�*,��*�d#��l*�
0BcИ�V+8*ϸs�.Y�QN ��s���}�޹�u E$3���[�wIV�%��.���k�R�&`P"�D�u�k��',�g)��=��2�C�6�(�H�R�,Ǟ{��(i��~l#G?��R��ہn��w�)]0��襱����w�)���|�� :�����]2�;�~��e�_ �n� :8q��&�gY"�њLD��VRZP�������~����O5��ڗʞ��T �S!2��ǰp]��9"@�D�Dۇl1S��6JK�.Q���j������*��_��W�
��3N����}����M�HZ��v��|�����Xmuõk�x���y�7�˓F��������c��%�n����#Ƥ��̍���_��Պ��������5�=�u]�컒rw�Qv<r�.d�>.��4��uY��(1���,�,��yX��e$��!��<Ϲ��Vg��9?Ƅ���1��Q�\;U[�shR���cd``!B�ȭ`��ߪT�Z��uR�h���!��A
��
-FC�IFÌ<�,����Yׁ:�[�����w-�sY?�ݧ�cAGr#�(�@+�tA)�'��I��̀I6b'+0Ab��AU	4o��!�E��C�%=7n� V�z��v�l�ݻ����v�"��[����/؝I� ��[[�����,D��� :3� ��(��ِ���ͦ�|!<�Gx��c+�O��g�����W_������������Z˝���|��I��u�ٽ��#�_A�֝�B�~���`$����2Fv&c|ԞԨ�<QD�V(�m�4!9��e��)v�'[��ܔw�������=w���q�6�J�-��u]?R����9u}E���("��>����Һ�r�J�bBD�1AX���ڷ~��|�G�	p��/|j_z�T��Jʳ��� �XDi�@o1(��l���2s1�25��o��h�n�pas��	�T�W�����~x��O��w��htH����]BsnJ��|�(��e�p�A��FG�"h�Ŝ�#j&X7��,����������c:9Z���j��ko�91X~�_���Q��|t��[�'�L�.{{���M>8�aS�L��`4(�Rt-k}�6_�R=z7���"��Is�����F��E�923    IDAT��a��}"S�3NΎp��DIUUH��T��\\t����b�ɠo��1k�f�b�YӬH)ט�>���]2� 	a�d�TPާ\����.;���+��L��>��3�R���f8,��&��K�JA-�2eHQ!U3 �į�d��k��פ.�4JR���Q��s��m���Q�^��Mb]pr�a�ƴ9c<�"c6?E��h4$<��8˚$#dMN&Z
��1��2)22�/���+��2�p���W��F��#��+��E݀@�0Z`�@���9�7w�B[�젅&�	�J�5-�Z"�Lu�~�Q�aA,-f�!W%�mL0����Ƃ*dM���iSsH����
�q���˺ϡ?�y��g������\Sw8�{��BF<BEv�y�+�\}v�`��w�l8b��ϲZrzr��{���w�ِ�%.�Zi�p�q���K��[����|t���������o~��vd�{��݆7n������Fh2�ϩ��9��x���P7'K��x������9 y�*L�b�W��jB�qYC�A,MI:qa���nQ��<UX|c�9�҄�D:�S��Aw�� X*��i!u]SU�:��֮��4Y!��1M�\hvی�D�w�k��U�v��#�������{}|_�XҳWkk-VX\+'���`�@{7'���$�r�L]=X�b0j��"E�Rx?�<��;����})�ɜ���2
DPA!�"&K
�պ��I,M� a�l�Ǘ��t~�B�X�ns������ZK�+T���d���]��%?��O0&��H�mp�rx��׾�7o^���!���|�������p��}����p�����l�6����stt�l�@J�.�Y���Ų�xmkC��z*�oG��Z��9���� �m�*�׻W�������E�:����-�~\y�m�AĔ5�ϧ����;>>��ÇX[���CYm03�g�����MfX�6��:|��V�*8B��hR��#ovM{��3'M�0���4y��ޟ��'L�Ӥmy� 	��᧿��B|�o-���1�=��2�����߈�����l;j#��<u��m�j���V�M��\[+�9E�>X琤�R�ܤ쉫+NOO�N���9�o�f>�o���,ţ|r_��`A& ����K���>���|�{�s��}��!U�� �@J����(P�	USR-�9;�����?��)�ߝn��ҟZW-rcȔ��Vܽ��Wy����وJ|��ort���`h��Z�)��1�N��he�-���˔�`������6ӿ[�- j�EB�J$JI�4D�xj���u��Z��mw㷿gte��-�\7�
�1$R��֦.�|���ϊ&�Ͷ3دh [N��t������0��	�bww�3V�eY󕯼��h,��yQ�Ri%�R���Nc=-���g�J�� Hݺ1����7��:�3�ݜ�v�g�  @)����i�dQ����Op��k�(<�/O��j�*�%�-�	$��>3��v��M�9�ވL 3� $쵀����i��������	����y?g-�p��#� M�`����F\I)���?�W�ݼ�c�蓎C����k+TU�{����ﰿ����s��9L}�� ����X�vv�������]�R�����C~��1<�X��˗Y]]mnސ�a�댛뺤(�MA����O.�>���	�/���S�p�9DS��pOR�}�c�puͤ��Z#��p���}PN/x��H����pt�ϣ��2���.����)i#�ik��*�ڢ�	B������nۻ�plx 
BZ�����5�W�:���h�r�lRQ��Cʲ����0����XWRW%Q��R�ѓ���<��K���O�8sp�ǃ���#u���6��IW�����Z]Bb]՝A������r���p#�p8D�U�4F��\< )Rx�18Sa���y��+�(�y���n�b>�#��T����.
?��צ��>d,Ǫm��£�D	��,���z������7^CĖ�9i�Y��*/*am�kCʣC޻�BL�B"�"J�$��V�ID?��#AY��{�%�b����q��W��M��O��n�٣�=J;"�P�#|P�.S�_��{���7��N4�*���I��c&�!*2�P��l-�鏮�]�+�څR�m�.|m���Сut���Ű�!�|A�9!�ɹӴ��/�n�Y�X,j[��ח���p���������`0�,k���)˒�����W�Z�����qB�}?��sc�'���O�������b�}9>����H�,f��%�ً�l����Xw[�H��^�BI8�� x��$	:ߐ	�#�5Rx����R�q���W^���+X[����-Y/�Ҷ<dooo׮��/�@��x��{{{L��N��-�89�t�C���5���Y���0n�m4�l�2���i��k'���,��l��$nM����i��^t�ߓ�	��{��ߦ�O9<�G)	ޒ�9�p̷~ɀ�!Hw���4�}C����Ǐ��ˊn�,�l<�p�5oj��`m�1%��Ԧ`:�������!��״���ԅk
��)�?a�M�ע}��������.yp����Ģ���7o������9���������
�Ǜ�� ,9:�FɈ^?�dIg��Dw�4��x��MP���Bx���.���oY]]����<xp?,^$S7�U���00�3¡U�	�]����h����Wōb�b|������|F9έd��t���s��w��}҉T1�%�T�\������B�����&/�>ZG��=�:bg�����l���y��"�s��%Dg�&>3�z�5�u5�G���Ѓ��Ak���ۚ<ː��L�@i��e{����Z'��_�)�_+<k�4M�� l�R!�h���0�
����d;cʲX\
-e����~Y��n��k����&�	���
����g�g��ё�L����F^:Q�z\:�+k�a�#�/�w���r�,�� ٠e���p�AVJ��ټ<e�Z��l4�[�;�B�׸z*�H�H��ш(�(˜$������������C66W���g���3�������e>�G�[��(��#����l�SI�0)k�t:�$�D�0[�Z[�ő\>:�ǡ��^J)ZT�S��|��Ok,�
=��]ݿ5B ![�k�̡4�������H�g�)2���Y_��=��pM"�r��^Gm�(B�A��£A�T�u֕8_amIY�p�0�g���P�9u-:�x��΢��8��찰[ �$/N�s�=<s5ݢ��t�Iӌ�h�$I������&:D#�GuH�1�4�H��a��h@��U[$Ƒj����>��t|�/���q�����	Y/���R�z)e�?��|�Z�
P1�&SY8��Ԥq��2�m�����X];ǅ�A���%���C2�IJ9?"�,YoH:ai�JŊ(�w�҂~��f�Dc*��7����(���7�@�����=��#���^��hfӊ�k{-�"���h%I҈HKr���(x�?	uW�H�k �"�_0l���4�n����Py!:ZBK%i3����5ݳc��l]Ҭ��)�<�\#fA�|l/�
���d7oE����@�mO2��������I�1�����a0��?�w���?�7�@J%�?U�����+�|GR�U�g�z�ϻ�����~r8焋��	�����^;V�=k�\�=����c1[.����v/�i�l
*�5����`D)f����cl�o��7��u�y�wl?z��!zK�0���!:R	���p|r�`�#Mz��c�8���Q�5EQ���z=&�IW��� Z�(Uw��{�@/�!�F<��(�$a}}���-z��P/�(._;�󷼂]F'Ϣ{�{�%;ۀ���t�a��q΄V��x	R;�ڰT�6+��O�kF�DhW.���]��7�� �X�\�?	�(_S�I<�U ��B8�j ʡ��69y1k��,���Y�5�O\��2H�(�)Yo�J"�bwߦv%��,�(jKE\�x�^x���M�$��
��ίG���H�\�t�˄βGH��)�����"��;��5E9eZ�C[Ζ� HQU�z>-B��#�'���k;6�'�
t�$��XW�d�d|�/~�S=�a��%ta�E�#._����\�r/"� �f��;h����R�,�x���'K&�}n�>J�X�or���Aµ�����(&������dDD$:
h��p���\Acp��eLxk�!�z��by��z�E�vQ�=+�m�s���R\�����ͭ�W�u�֓$a���Ÿ)�H�p��.z��M{��\ӑpg�ݟ�tY�sJ);���xZ)�9:<A*����ß�ٿ���&k�k8�y����|�����y.�2�x\���NƫZ��*��y/�/�{<�cC�$�H�{�Cs������ܾw�\�]}T;����27�)���KE����4���b��d��T3F�>[�׈#���ڵ+�e���;�*��K�$I@h��G'Gd��,���$I�|̙#�t�܎%��
MܗpMK���-��$���b�z=��{KQ��,�����E���#}X[���^z��Wd�\5��%΅8*c�MF����~��qO/<��+A����f�ǟ�N!��E�bm��AZ����Y%]�^`�����Bx��g,x���Z���эi�j�oQ!@i�w5:��y>�xC��A`a<�~�˗�r��u��~��*��)��y��:!�����9�PQD�#Ԓ�H)�ܕM��7|)C0��iLU��"CHRTd��ȃMt�/,Z��s��N����炝H/I�.��zNGr��o�����h��G�$��`��/��*?����À&'}t���T�Li��V�R�,���S	�e6�p��ۤ����&�%��fl��1�%L��G������;4�}S<c �|>�4��`d�MXT�3���`��8��>��ܙ4����	�'�
��3�罳�-����P����8f���M]��g���B�ݽp:�m�����p����$�e����U�慗^������޿����E����l����'T�%k�ON���f�p��o���ّ���������8�� ���|B|\����y��&�m��l�p
-�
0��:�o':J��)5ei��=�ш^���ã=�6���~HQ�Y]q|b�N�E�x|�(.�
{>�vm���SJ��=��RW�i1ĝ�_�<�b1�ڬ-�<�ǎA�HR,��Hwj�e��PB�z^���/�����f���l�c���
(h�w�E��ؐ�!�,P+�v#�@���x� �g�>�pq�R�A�~4�_���_��x����	��U���(=B��Ƙ
c+�(%I�"�����-U��-G�$�X<��^�|6�Z�"M��DQ��|�#U�4MYYY�r�[^T���yM��*�D��'ME	TEG�B@)��u�#��7� )ΦAJ�Ғ���Ee1u]1�N��dYFU5|�S��pm�?�L��o�z�	��H�{=I#tB:��b�!N��g)�����c�jfv(���o�k��X[���
��#Bb�R�q!=RA�UH7�X�� ),G����M�^����*����Wz��x�T�y�uQhѱ<ϙN��u�Vqb�Ž�H��w���{\�pCגn��)��Ej
��s�2��}m0X�\b�����9��.E�U�.[��������i��M�|ip�m�T�<���SǱJ��������o��K/����XҊ���ƍ�z=����r�
����]�u]+))CI���[�[o��%��/d<W�W�W"�8a�qRD�*�,�cP���^�����G�u]s��e��~C`?�����4M?���J��O���2qj=#QAҴ�wtF
�����]h��Q�h4"N4U9�~�cv�k�����~IQ�qƲ��M�Fx'������3��9���\<�۷owh��񄕕������_kݥ3�E_Pg��7��9ٴ��ޓei�bmN�)t-;��0!'���!�x����*&�6���>��g.�s�>lϣo#�AW�5)*єEN&EG�|��V��!��w U��-�=���H���a4�ĺ�JP�K����>\���eN�X[gZ�@QU5UU�kT,�O�j���>�R�����.r"E����Ue���e�
��������}�����+_y9�9ͥ����
��/��n�]��BX`���c��L���2����3T��~kmC���������X�<���a�W�K�ʃWbʺ�zE������c�X��:!JRfSà��&�	i��%	��q8�^�kV��^3�`��]+e���eN:L��qrN/Yc��}���?!����_�7ڢ�'�B1�b��.8hqc
�kx�H9VVW�(�g�4^�?R�4ee�����:�'3��)�+����g�Bт�!�[�����,K⸇֊�*O)w�E�֚���Ά(̹a^L���ڊ%���`0 `41��-W��W�!�i0���NY���c�$ass�[�lnn�2ڠ,K�޽K�$lmm���#��9�� �����ϟ���<�y����w����Ue:�<����>��6�����R3��.���(k!���j\��[o�u�c�_�/��x1l��.rRJ��!��{!�Ctj�g=����p���*eYvR�4�U��SѐjC=�lo��@D][��7d}}��QG���G��,u]��:
�#��xb��H�&��7����t��YAQZ���7���[ᵫ̎ /%R��Izy���B���e�}k�ܒ����/�h;v�N�[~�?No'�4MI���F9�������v�פ���@h�FQ�Pck�
��BL)�����q���C���gg��'���/֗9o��k�����V.��p|<���)%�Y�|>'�Ť:�,g�\�φ�c��*7�%*��%���.�э��sM1�	|�Ó�o��,��g8Ҵ�Z�"beu��h��|ʠ��7G���(퉵���3�X����h-�g'���?��0�!R��Sa=�C$<�/r��98xȍ7�<_ya�A�`�D��Q��	��#/
��#/B������67���!/K�
��F*�$UQT��{�a4X�_��&�^�m���t����;�YƬ�hP��e��cNM+��L����;w�<\����j�vk���v�P*�R������0Y���z�M��������
��x̵k�XYY����{��Q_�����׿NY�ܽ�����,���{ܾ}��lֵ��c�w�9��\8�R�ⱃ���g=>��#����(�9'�t���>�Z�\~��ڶ��<���ڂ�I\��c�p=��cyH/�v`}/jՎ�l�����q��9VW *lUr��<�WPy@��-�4%�"VWG� s6�6��v����z����!�������X�"��-a�Cv\k	�ϬtR*�q��vZ�;��v��E���,ӳZ��X����+�jS+I�$D͝`�A���l��V�'��h�Pm��2V�p�!N���uЃ7�0��]-#�tqv>��}�t�d�?��%%��-m��f���6�Xou��s@���&��3��L��j�v�U��B(�X��u
![���"�T��M|��Zy�%���p&��,�B�H�n#�~�CE�աɋ�8θp�*k�[���*
����
c
L='�)�������_{�e���]��<P�Q@[#�p8R*��J�DxI"�ق�b�g>+y����%��ӿ~!�H��TL*��(ͨJͬ�QQD�E(o�r�:_{�޽q���Cjc���'%�� qD����~�+|���y��5����c�ݽ�/�s�ܹ��GO?�˭�v�߷T��(�⮋����K�\өq�u}rr�xr@�e"�)q�q��Z�|>i�C�1��x���Q������p���z�%;��Zs��9��kkkݜ����ŋy�׸t���ܥ�-k̋P�~��_%���w�yYS[h+:�Ҍ��Ka��3!�!����e������+��@��{JJ�Fz�!�    IDAT�{�kZh�����c��<�>eY�]��J�i� ���>
^bNڮ���dx#�d逵�67G�R��!�uf2p����F��3�i����e}�!i�����pttDY�$IF�$Ե�"�Zr��-Ue����C��Xۺ;�SEA�&��hbA\>Mv���RH6"�� g�zZ�x��
=����E9 �M)�w�)�C[�k�@�7ކ�)��)���v��E�v��:�v��`Q�dԠ{B@��=X���<u(���R���EԡގP.�S3 䂪�Y_�`}e��ׯ�#RM��!�7{ё�E���+�ٴ�'d(R�u�s`}�ݮ��6"�.�~���"k+*Sb�'�R�b���׿�������g�lz�|>�N�x�E���	�ϭ��g|�O@I&������ܹs'x�	���x�w
SC�N*� c+�g�d�`�;�X6��Ylr~m�ee�ޅ�T��NҌ�L�����4����.���}����<z�<�69��A���k���:���&�뛬�mP�5E1gw������?�1�*B������D��A5)0����ϝ�E�ϟ�d�t:%�SVWW��stt�TS;t$I�^��
 ��1�O(�^�h�JU$qF�FL'��N����s��9^x�&�	{{{L�S�1dY��/��w���R����|pg��/�e�yAkVVV��w�y��n9�a��B΄RR���������������/d<�zw�Z���.Fh'b�E)^
�&����1g�7�2����jUP�;���YV�N����>���.L���*[[�����)�6�p�2�M����	�X�,�ܔ
7[QT�e��G���<x��������'�s�$aee)%��PH���[�!���W�D����}ʘ:���E\���!t��8�����X�7y���BȝQ�6�^�cl~_iI�e�#}(V��(a2�
'�Kdѫ`� !��#}c�,�`�9����ؠ�E"t��-Ri��o��A�#E���g�������O<�X6ŞpOR���"HVV���7�䅫W��S�,[��pO�:�d�T����ĲD��
)u���'�"�~�l��l8�A�{����F�1��i6o���ˊ�����]�_;��)��/w���<|p����S��#��6YY���7�/}�Ud/a:=$M��}�������Q�BH��Y0zd��R�%��	�	�h����1DB�瞻w-�l�Qo����YJiJF�b��T���jDl1N�Im=�2�G+���-._�y�c�y>&���qJ6�&}��h���j
��>�����׼��;��:j���S5��Bt
�6�m���pQ��-�~���z!TJS��$I1��(Jf�)�露���{TU�����\c�CɈ��sD��L�ۖ|��Qy�wԓ6`8���	��.{��
R�e��W(���7o��H���q��^�=
!��H%Ơ��
����2���k���DJh�X0�}��]��=�}�����$鐦��i��5>i{7�nИw����H��b��367.p��UVeuL]嬯�S����f�&����Ƶ=�1��U�(q3�����`g��,���*���7��q�"[v�7�4��c�E����/��j�Ek��i(w�vN>��h��U6��SzM�P.dAl!���@��+�� �B����}ֻ��N_*B[�
"I,.\���9�R!�-w%q"�����k}#
���e��G�!�
���]?�}�g7�yE����˺�Ը\2��ڵk|�+�p��y�j�mK8��L��k�m��k��N�nz���m��YxHʈU�E�DIL�H�>�����E�aHe9�������W.l���`�5׮_a2�g:>�*J��D:c�_ޡ�����X�(�G���������h)0U��B��t:�,k�h~�d<g���$JgX#��!��~�w��Z��n�z���&�����u�ԜL��Uh#��"d
u����c�pD:ec}�nUR�S0A|��2��r2�b�GE1eY����O~�c~���SU����i��\���e��5a.˒�|��w��҂{mm�_|��xʝ;w ������A�M��$I�1O��ʾ(J�
?��666�R0��h��x����8fss�8�I8��=���tH�ݻG�\�~�<��ƍܸq��vm�]���1���766��o��eǿ��\E_m���v�:@�@�RI�r"���=�[H����8[�곎���}��]�:�eMU��<��y��@r|R3��p�,;�����\�r���5��)���[��r�w��9���ܽ����}N��R��X]]Ek���.'''$I�e����J4����*���->����=^���O>���w�����+�˿п����Z�F:�
�X(�������</B�֫���@4�7G@��V�L��;�s{f�p�$����*��ƣ�`�ӝ�%.��is�������Q# ��g48T����
_׃��3�c{{�|:Ai�|�\W�i)�.X	}�l���i�K�M^P�j!���DЅ'1^���ț�v��SCu�g���w皮m�O]��p�&/����?o�ƛ�s���m���>���Ջ\ؼB��ump6(r��)�uă!��~����o�����G��\;�xf�`:�3�嘍!�d{g��}��T��e���H��*���)^&��7޻��`�H������?���gQ�B+*�8>s��
Q�����xj�+�tD�`�lBR;�`o�����;��m���YY��e�uIU���no��`��v�B78O���H��TY�M'�/��� �K���8Nq�5�^AQ,l��:�&M-i1:+�V���y�3l�ᬵ$I�����C��@����=N�˂��u�(���9�Yjk�D�&;�3k;E��я���S�������H�sBi/�PBJi�.<8E�mbiE���K)�!b��z�4-s,�g<O{7��<�D���;�,KI{0��u�����F}�^�ʵ�3�N�˒���]8O������׿�-{G�$�ek뛬��1��893�Y[�h���[�Y���K�e�/�B[�"2/P�Ӧ��b!��=�����}�Gl=�
��m�h��"؄���{iz�$�eKhLӚ�h�q(!2�x�bmMU�H)�W��s�7�7m��\�E݈�G�%�?�aX�-��|Z���'��%tԇeN���oݺ���#�8��s��Y�^T�Y�	�7�\
%�:>p`A
�p ��&Dg)�2'�ׇ֤i�S�e�d2�,�ywjۄ�r��4�-P"�ރ�TE����M���6FԦ+��xop�RW)��u�DhE]��������.����gS�xE�:ؓEX8V���CƓ�y�P8g"�������W��[>�����VV�ܾͭ[��̦H����3�Lx�h�������T6�c#"G��CV��,��	4��䓒[�n������?�Z���j�zm�"$������{�庵ܷ�a�h��s�$a6����o�����$	�����j���eMk��q�z�eeYrtt�|>��_�Z�I�0:�s2�t����ۦ�lmmq2S�y�w:88`ww�?��?������g?����.���B:�]�p+�l��/�?���E_m�L����9Q�8V�>ʍ���F��DG�<�i�cpQ�	��e����`�P���sDh�Z'I�U���N#�	 Q*A�cBJ���j����Rtxd8�_^�M��y�wv�ȁ���d����ܻY��"�J�[�_cw�psJ��q�ҋ\�t�G0�?�dg����M67C+���ܻw#������k��1�s|r���Z��"�S�ӥ��S��Y�m�kreCFr�1P�_���&Uh[C�C��d�MVd��|H}BӋe��Z1O+��OA� C&��|�><yq��ƺ���I< R�T�GD�,`j��b�^�#6�]ccm�)��cU��4R%���c�$l�X!B¡���%�[ba�eN9�G�>��H�^<'�%B���S(J!�¢�EKA�<G'cD�%C&�l0D�����-�Z��Y�׶ЯT�����H�P��v�pB`e�P���H!Hc�)r�|LgX;d|,�	����9��l���A����`��B� pr"B�^���+����r�zN;FIƴ8��H�r�2#B \N,���)uY���^�э�Z���M��'�~�uQz���s�QMP�` $��}~��cNv��Ͼ�o~����$!���%Η8�k�7�y������_���Q��}�V�z�kN�czf��dʃ_�7���g?��ܕ�B��З�K�Jcs�4�H� I2�x�w���=���>'''�'B@�G_D������� �qK7�AtH���:�^Hp1r�����#}�-��`��&ZW7�8,��eG�,I�P� ���ׂ���4�ac�!<��
Q�'Ix%��$�Mf�	u=��_AG�a6-H� ��)�+�p
8B��`�'�F+8�u����35�Tp�Σ�$f6�09�Q"���P�N&��"�bp���\8w��sx`0u J��yI�qIQ3!R#�Y�)2� E��;?N�'�5����_���я~�I�޿_���E_��;m�y!�x�W�[��y��Y��
�۟����a}-��JRX�����w��������"J��C�:��k�X0�������Ehlmm�ꫯrt����i�t:����loo3���hD�$lll0��L&݃��W��z���e,�-O0�?�W��/H{����AkL0�n=c���X��$���U.]�ĵ+�Q*ؑ@���������{�j⤼k�=��FKh�0u@�A%8')�c<eY!�"K��C����A7f-�8d��U�)���p��s�a��G�P ��� u
T"I����Hc� �h�k(~]��@zZO@���X,"�'�8L���ru�{�N��ZŌ�#և#�sN�w(�YE�k󳞌�2�rHx�Rz�j��;7����o8�"Q�%���5Ζ�C*�������������%����Uf�O��O�͛�(����n_�����K�c�R�RAY8�u�S圌UY�_��� ?���
\�5v�D�T�M��+���Ռ�*��>)^��-Fh�6�[�:�D* �
�-��V�I�`�
g�BL�1E9�*U]�l�=)4Λ`g�O;�V��F���c�ܹ�p8ll^���
NNN8::��իH	q��c�ֲ�xo�L���P�U������Z�S����0���oZ�WF�QE�M��':�_�/�x��#��JL�ｗކ�+*��v�mզOg�C�k�i]z�rw�Σ�Y*�"�x|���3���ˬ��o\��>��`u��x��ct�cw����;��Q�
V���[k+\�|���-�s������n��޶��� ��a5ݴ!����=�W�l�v�ǭU���j	���������b#L�j����A4-��[H8O��|d����ۺ���E9���T�	�m�k
i��Y[nՋ�M��R�(�J!��?0���d���>��P�B���I��R�$��X�	�����I�/]��ڧ޼gc�����6�]�h���A4���*1¢��a�����@^�������2�8��
��"��rw�*X4"��� \�
!BKLـ�{B��V!��Mr����{���/��M�^��)����ȝ�ߡ͚������O�̇+��"dDGo���|p��7�)BJ�g���]���������h�XOY�sgkL-�#�3��wnq�w�Z�e}�S���J$D�	�����{�K�8�RD*9��Ԧ��΃@u����A�-=�m�89��!�2�V��'�^�w��8��K��ҋ(5U�1�ƒ	kPJ൦��࣮J�8B)��hN][��5��'��TU�3��P��JE�klm�u�q5���AG�Z��f2ws����$x���EenQ2�ʕ+!�c���l�e��r>X"9�!�C)���D����U�EZ{]
YW��*�s���e�VE���3��\��{v���HN�"M���������o8?�����V�׸�R
Q�������.��qtt�W(-��bv�<���f3����`����k�G�8�"��޽��Qh�dY����Y�[O"з����;����4?��?a�Ҏ�3RH)�|������;���>B�< �q�R�5'�)�*q�P�-n�D	2��Ea��z��������=�$j+�k�����}*k�+�s0诒d}��*np��j7$SHLT�E�fߟr���=,l~�X2�>���$�)�Z���DR!��U5UQa�G�4��p��iS�36l�w8b�p�" *a��8A"p$�uH,J���օbNhjkR��y�7���]���g�c��e:>��WDk��Z�|N�,C�Z�6�u�,�����!&��:��U𜌢Z�]�0t�`"��KZ�4E�R��Q�,�b�>j��Z��mv���Jΰ��ƹ(�J)��!�E��`	~�����2�rh���P�8��0��\й,<�8�i�"�u��WW��RjSrr�d@7��$�J"EP𛺤ȃ�6�����c����4~�g=:RX[c]��H5�3�XF8�I�OӔ��5z���T���u�]�v�S��(�Nk�ׯ_g8\��������ˠ_�sNHD^?r�?���s��]�_�/��X1lxo����ށw8����[ŧ���0�^����mW�4��n����$Iё�*s�}��e��䐣������>�"1V����!��`����d�ݻ����X���#N���'�F�΋��r�����{97��� �g�E���S/4K�x�����޷��l|��llm���m6�%�f��W�d2~�Vo]�����1��cY�eY6�����lk�[/qޅD����N�m^�0�����9�{�N(+H��N1UAU���\Y?���*[�xW1�3�}�No,^�<�gi�x����Q9��:���$�ܮ]�ֹu^z�%F�!�*�{���7?@��Jǚ4ӤYL�hL�֠T[ny�M�ƅ��&� pE��;�u��!����|�B�Ƃ�2���X#�2���Ο?O����p�i�R=��S���G�C[�Ra���!�$R1+�Оs�x���\ݕ���uU��yn�nh���K���y������siKyP�1�k$�������Q,��L`G�"�r�k?$�!d#l*�X��R;��}�rY`���8g�Lf8<Q��T���4�#޷Tp�P�s�*u�J~��!�Bk�X1�0Gp��a��$q���.%G���tʅ�h�%�akѴ�ei���̦ަln��_&�2���!�E/�{����[�ȸ:��ϻZ���i��U�E�H�z|����g5�nˈXˇ;��O�֗T�H��)�Ȉ(N0u��7GQNy��>��y�/����pm���&��)����bw�$�$qȷ}�hֲ�x��js�����c�ݻ���4Mê�1m�ܜsO}�/?��|Z�H_;�{��EkW�9����u6ϥ>dg�7n|Н�`$l���T��1e���æ�rݤi��p��o4^�vUz�ex��B{L%D� �$q�f��H1B
� "�z��mq��6�G�ń��-D���AC�5*8k��c���<]|�����PT�._y���/����&��	o���<|EN]�И����*��d$֡ �B�����(��Ix0��z���Fk����2��`�(����VV�HӬSOJ�9],|�����є�ߴd֖�F0�.����f�u�>ȶI�-EE�s���R���˧�r=��tu���,��B��s8�R^��HJ���=PJSzYڨ���D�t$��l�1�,]�U�aU��Z�bzα<��=,
��p�J���$�2�@�8jP��؎"��I�9�Y&��2���P�7]&Ѫ���P���2M�\eQ���O�����    IDAT���Ԇ�BE�^�Q[��d�ݣ�h���!�-�s�����k���sOe�ɋ���Do>�˷�*y�u�����������]�IQ����E-�wz7�`]&�����~]V.�����KHIk8�M)!����	�]o=BJ��y���7���ܿ��/_�W^�ҕk�C�
�#�*��!!�Uak��d��考�Cd�:i=[ې�����8>>fuu��ܵ(�2b����Z����(X��I�0���9�Ej���H����[��j泄,��d_ꪤ2QST+�dY��/6~��T�Y��l<�hb�N�f�=�I����� �Y�G�*�:�?����tF�KA:<c����8PY��4Ր̽���3�_�-{�M��i�D�pT��NJk��u.\�ʅ�5�Iƃ�:�����fK�$Ǚ�f��g�%#"�2kA
A�
��閙���6#-���as(�&� X���K�q_�L��������\�P�����Wsw35�_��T�zEJ�k���8=;f<��i	;��%�=$&��F�L!���Llq�������e8��*\�K�
��z��(�uU�F�����Fߎh_��!MB3g��"c�R�&��_��s�h��$�H��_Wh��z9�i%ƾ� ��s�#��T��wl�*Ꝺ6�i|`��o8}���"6-o�M�GB�zs����(W�}���ZKD8x�o��ggԭ�e%#14Ik7J[����A����F4��$;^�������%��7�&R/J�+�TiL��{�0�r�F�F�	�˪�����j8xu����'��ƛ��h}��MRoÙ���b58������E��_����gj�k���sE���q�j��TDt8��CY�޽�_�1I�(�0 ��]���Ʉ"MS�J��Ņ�('g�{p�������aww��tJhjvv��7Xq�JY��'�X��O��h8::�6nݺ�b����:mF����6F��1}���Ί��<}�^��8ŤX��R���p���,+R�C]z�y���6k�5,b��?ˌMчˑR1���0����!�u]����x�99=b�\�\�h���^)kOU���h4aR�t�4��Q�'��WH�iGμ��6J\>Ƹ���>��Yk�rK�;��cLPW�D/��5!:GU��Fr���O�0*uS��y�&���ɹ���Ȓ²�9==��|I�-(AK�۩"dYF�4����K�}{�y6Zs���3X�D^"aP�Fw[qb#�"�C$��/�����|>���ʑ�%������R��鴏���$����1�k�HB���Ɛ���7�xc��Iz�I*� �@Q��k]�Ջ�U��a1G1��������O[����.i�����3�l�b��Nz�Q+����ELr�TB��E��X�{^�=�T�D�\�9˻�ڐ8B��>��!G�f +�x��o��?����ۿ�?���NE6u ���0���$����A�AU��9�I<��ݻ߾P��}-�LN��i�&�� 0b��(���0�M� mp�O�1��*:C����buI�n̼��X�sB�r)�wi0%�UD��-�FŚX.�X�	wr>������L&�f3��������H�h�4�r1g�8g�� ��Î�S���y�Z=ٻ�`�&��S���v1����]���C�`�4��q��}����/_����p��o��S�l������*�������w��DQ�u:�&b�a{{���{���?����px�"˱VX�k�Rb`�Z��Y�	��-f)u��Q�Ν�����VG�"�G5R�%*�&6�U�x:��+><���o0��&����������K��xL�˧}���N"��I�[5/�u�|4�mEȲ�,P9�3n��g~�Bb�Ν�L�...cs��f�Z`D��g���E���)�#vw����,��`�Y�
����`�� ks�/P��1_&�k-����] &�IOXH��*��ϵ�0s�>�<�=�z����8��2x!� ����E&[�lmj����`u���צ������z�]thX�}'ǚ���.=�>$bmR��\F/��ϡS万`��@�o"�vi��:��E3���];_v⾲y��V7u�s4u�K���S�����O�ۿɽ{��w�GY,E���9e]��#�|����;;ЄN^-I�9�R� e���pĨm�Vڬ�e���ֶ���_ݥ��I~j{�K�mmm1�88�K��0�Z-�:�A��՝|�Q�8�IفT�8	�ߔ��������m�?\��bϞ�5Fc��IPE��FU�����d}q��i��j��{?,T��cJO �����b�����|b�O��\-�,P]2���h\���2�,'�i�1�TAhj|]��e"X�����^F!E�5k��!fo���9��2�1|ݘ���y��H��6�(��qy��M�����> y��U���S>��C�5�Q�%��Q戡�)rG�Y|������c3�s9M8??������Z椴Ѡ--I�T'�:u�J�g	[�����1�0�&�'pn\akmH�s��6��1���S��Ӫi����݄�\�-�g��}dk���[��1r���w?z�Ç��u���� ��˳�^�&'��� ���򐲊�z�~rNc�����*ߪ��~�"��h����E���37�T=����>'��~��V����Sr�t�o3z9Z�QP]a�z���?���7�q�Ǿ����Z��^u�_�UU��kqy�G��>�{�d#v�n2۾�[o�`]��~��_qrz�[o����{+�R��I���J}�&����4Ep���R��)�g-�ṷ���2��s�dY����܄
�2�)�O���d��D6���,��C��*D�چ?�{��o_}�����}��Y��Aϐ���i"Ĩ���vn��:���U��u8�LY�E�J�YBS��K5m�.����^�ΰۊ5��MZ�t+-'�q�Ybh�c:�my�4z,I��� U"�敽�#��(�X!AlZ�s��鰜���fD�e�����ڶa3�U�b��5'ƥjHqX��E0Zy\"��N!rz��s���ɸH��1�!�����Ua<����$��hR��������YT�Ծ�	5j�@����l�ɇ�)�kmJ���{@c-�Cr؞ކ�޿���m�5���|�bQc�8�������F
5�"�$��S��)'G'���;����T�yn������	���&�-b��V+Bp6�(�LFc\fPm���Ū�,kn��:ǯ�����T8m�g�=JQ�֑e0�ʠ�;�*�r=m�^���������Ē��6�k���y�?�%�9���_e��ĸv´K�>����f��G�߯/-���I�Ŏ*�Q{1�/�s.�	-ԧ���tZP;y�""qMk4�VLg����������&U+��	�4MCY�}֤s�D��h�!/:�t�eh�����,F,��͕�o��:�ҝ��c�*���g-�Q��朝�%�WǛ�T�*A|1��h�yc�v9���GGx��}#�\�>1�bLH��h�4���u������������t��~�����j��N����z �1��)�D?�^h�bM��9�X��7�/���:�V�t�&�ۑ@;�в��g|F��q��k��"��k,�,�9����(OSG���]�G�<��6Q7t���Ʉ��m��xRP. ʍ�=�g��i|�3��nN��'�
ʺ��!�Fd�4�ȊU����prVS5���і3�f�,s��`]�E%�{n��i��^��N���t�~
-���g��^�|�^�=E�k�8g:�2�LZ'�����rNӔT�_'���l���=f�m���lIU՜��pq���R���D�!��4�r�����������X��Y�-��ç>z��iˡC��1v�i���4���9|O�0�����A�n�fi�2�}������`K�Mj������u��f�����Nx�i����K�/fݤ�j1�ĸ�uϲ�Xe�8$��$Bu����+.3�
��F�]�nȍ0�nq�`��I)z��ɰ�`�����6��7i;��Ј0�'};w�u�	x��|_�d	���9182;�����������{rxx���uT��i�U��\��D�ЪV�������1a_�wƞ��+K(\��[pѪS�(�����M���a<O��*:|"����%�*Gz��cl�N�`p�]H�U��~9�`�z]UM4�1U;~@Y�pN/��_�:g�q���'���w>��F��j@H���
�s�b��T>2��:�@Gm�e��J*.���`gk�ӣcV��q��֘���"����HSVI�c�3*�c�mHU��boo��(�ǣ��D9:>��	H����s����F�[�Qf[�:���u���dY{�����(�:�W���6a`��1W��l|�*���o���os��>��}��Pΰ�����;�ܿI����9��X��Y.眜�2�� ��l<b2as����a1_�������8:>e4�0�n���o�Z��֭���)׍��#�tU�=M�^��I�E�L���c#��'miQX/�X����:F��=à]_��+W�b6+�t��^/���c����\2B i|���`����j����A�n�~�����9��sv����C��n���K���9;;�В�'j�%�D���y��S���o3AI���x�����4M_`ש/ucbwm��L�˅�.���S���|ʃ���J�7����W�"j����y��7�J����1}"��N_�@�c�&��VET:2��e�(��һ�s��%�rլ�{��,6�;�iYόe8��n�?��4mg�!jr��t�i�:�����d��aV���_Ԇ�Ʈ��v�P.��e��y�q��E�����m+}2$"!�7��y�=�2�7�N4���<��s^y啄��}�|�5����8?9�p�î�|<��<�f�&����ck�1*�����4JR���l�b^��H&�c����2�Hd�loo3���&T�S̏s�z\g10m;��t?k�d� &�����c"pzzʧ�~ʍ�XqL�[��H��튐�U��PWy>�(<���V�"�!2�looc2a�UY�������>����nJ��bLh��q�i�ez#M�m3T,b��ω����˟�*R�FV�z��KP7h7һO�Fq��W����ٝWM�0x��� �@@/E��	������7M�#p��=�������������G4��r�r��^���s�>���N�_������HQ��������`B�������h����C��`��Y��������u����KwOuϠ�TU�0��+�DL�2޻q���%�M$��Tc�Ce$~*�֫�m_T�Jl*�,N_zG �[�jT-TԈؐ�k'�_�+һ_��=�#g"������Lb���iA������1��i���V�4����`Z�!��EZ�-�i$l+<����Cl;��s�i<�����0�ڞ�:Ƙc_Rvx]_�6a�ԆЦA5�DIn������GTָ�>�m�:ӟ�l6��A?�����W8#_R��0Z㌧Y�m����R�:��l�+�^��믃��?���^P�D�z|r�r���"��S�RMkgyb��s�a�x;��)n��9~�hf��ެ�E�,IJ'�iSD��'Y�UUE��d�`>_��_��������wf4��������8�Q�5�ɹ�w�����IJu`~v���G�D��Ŋ���G4��9��>�7�S:,T�Oc\b;��m`�b��^�]֞'�M��TXs�B?�4�}`�Tn�E����v�-o��"�_y�p��uI#>B�4�����e��@ދ�]�c�i����c.V+2W���~�F-gN�4�[5%#�|4�����ƍ�N[g�:N&#)-��#������>h"�6.��Y��ݏè�p��uR��Q��k){Ʋi��9F���};�Y�*ĸ2bVx]a`|�c
.^����;c�髍ё�ob�@FD4���}O���������s�����e[�aL�'��֮HumD�����������P�
=ۼD�>�m�vm��k��6gb/���0�������P�4���q�����4D|c͢�^�$ ��x��J&����{<M�e����9�W?�Ï>����������-vvvx���.W������!���Lfۨ"�\�|������Sמ��)}�^��1;�3�����6\RGY.�V���b���?�=.�$�!���u�,��t���	=�1����jU�8��jŗw��T%��2��5��[os���+|��(V�U?�؞mQd#&ň��4e���!�G'����Z��1�ęƦ�����W������v����Y�y�a���!�}��9{�J'":`���G5tYߒn��#�L�١|d�+�y�o�X�c>��'�(���N��F\{���ØV�CM��� &K�٘�2�/�X!�`4�����KCţ˰c>���.Ҽ.�3���1}�҆�	�����᲌�Y�Tvs����JU��>��\.�hGp�����39}۾�y�b�oauo��is��MY1N3�^�G2I��I�H�>���(O��^N�_��i�Ä́(�j��s@]=���YF>m��2�3���A�e��TU�)��G�Sƹ��(�\O�k"RU����]w�Wo�}��0v��h�����Rc���]�mM�*�q�MlFn�(7h\����qt�«#�r|P�
�qN�8����Ҁb��U���~�����U����|A�q�:6�9yh�����{_B11Gp�Lw���8qT͈�S��E�qc���?d<��ζ�|�޻���T��?���l���>O�ٚ�(k����(˒y]�}s�7f7���+|���|��g���<�����u������P�S�m�'_��ݏ���)u��{�����l�'���Ԉ����`" S�QĸD�'%�ɩM���9���޾�b^bl����P����)�{�67��g���/������?��r����9���|��f�n�����C&���~��� 	�b���Bye�&Lw0�Ġ��^��j�B�*�Dm5E�::������r{=-��I����Ϛ�j����^���a�4��t�|�
�[�/ɰhm��z����N� ������e7�=1�Ք8M�\r�6�Ԛ.sqUA1Q圭��O��l�E�N!\{���؀����Q��^i��
W�+B�&5��(+��?<Y�c���5�pb�pNaGԥ�.V�Te�J�d�f�pqv�a;֋Cʪ5�D�����m9�wo��G��[i���5�^����0�Ƭb�=Lt"��J`�R:�k8r �MD�W�� &�J'������*��)�#9E��m8| (HletB�rhq��I��E |�  ��vM8A��)nI�Gy֓z&,b@0D ��(1᪌ &i������t�0*����JN�>�ͷ朊}��w͆�䄏[߇]Z$qߥAŵ*[[[�����l6��4�����bӓ$�q��9�����e@r���{�������^����o����O(lRI0��j����N���M���/�h�hS|3��}?�N���_������6�޾�̓vv��~倽�'''|�ŗ	�8��n���::�)�^�L�4�#��B�A�}*ˈ`�
�v�=�ھ~�\�z9��}?|���~/;+�����q��5|i����-��>F%S�L�#b�)3�\,��ݴg'g�&�Q�h8#���D����3�` I��|҃+(H���Hh�Xc��Φ�G���9�˨����YKh&Wo�}v̀k�c�f��+�0��.5\.�]
$E�������FWfɚT�P�+�8�ڀq	�d�������,P��'N��4Q�t��N�a��x�R��� �Ι��ޣ��d�P�ȇ�����{�p��~+]癴�xu�`2\6�co͸u�^y�������{�����!�}�E��N
��d&�t��A�d�_�>:,n�/��۫R�y��4�b����=��o���%�A�    IDAT�G���p_WM>��3���|�rV�
I�Ay�X��Y҇c,J��'z��
^\��4MC�U����5a�|�_5x���=jCR���>+uyu����w�L������=iR2<����{�o�IOAT�(�QSˊ�k8�k�6�3;}���L'"���1���RŘˎP7x<�����FD#N��ƚ�K$4X�����W5�b���V5h��J���	K2_��^��^ds�VZ|��B�k��+�S�;B�QR䍎�?����l�����Z���@�^��f��"3�Pb�a�[vg�>��9��S�~�Ï_!�s'�A���I���X��>˲��t�R���;��w~����6�u�i�b�[Lc�m��@S�d�e������������*�5Tu�u��M��0}�M8�C�[z?�DIҜ�>6k-2��8�kO]�,�Kʲd:M����ϗw?㓏���Ç�:`M�1	C:_.����h4��H��D1��SʦS'H�^>j�V}t�9m��c�������t�ۢH��j�(��0E����U��{��l�yl����R�o8��!h1�%� ��K��|L���]�g����hM.Q� b�1�1��nVI¦ӇHO.��fEQ"F����$j�5cHd�⒟��ӈ�R���*�}�>� ݂t7_��&>f��!JΡ F����I_,�JJ��$�ISVT���D7@��`���|JrGѐecn����ɛo�f6��fNS��f�Gºk��~7��4�fg�~���rJ�k�,�h|�Ӕι6�k������.��$1��NP]y@�l����F#[d�A ��
[����N'hU�%�O�'F�?'���o��c$�L�d��9*�pZ$U�Z���>������!��Ox���s��O����9>�G�elMv��a$'�G,V�t����,<h��BL�Fg����X0$^�.�����3d��{�����[�Ӕ]�y��e{������w�.ߟ:p���w��o���Qc���(��]۟�=���C'Nѐa�c��D�-��qc�ߤ"O�{rz��qs�i��C�$��a4���
���k�T$K`n�o`�.W j���ҿ�H_��cΣ��7!`���S1��	m�"�fkUi��#bɊ��h��%,"4gyR/(Ya0�`3G�a���o��7�џ��;��Qk
g�)���y��6�B�v��"��6#˛i��:w���܍I������Z��f��k�1�N�Ӕ5>(��+O��XuT���sm1����6������՜�B�S�f������d�5��R��H�_�e����$|��]V����|���x��Œ�������������x�>xL���Y1����y���̗+���4��ڂ0�ku3�Dvxͧi�+qQ��k���cCxA��x�^^���Q���?��5���%e-�2�#}i���@B�^5�уj��\|u=ε���swf��(15��*�ڑ��Y���t�?顈��T��;ru4
�1�jػ�*?��@l��قH�1��󞾤�4��Z1<��?�B��.��jO�����)�ټd6�����t:m9���窍��F#f���,��w44�).7��#C>ʰy��##f�}�|L^�	V�
k���l+��%L�Ӷ���6ښuz�����ue���c %���)���0Ѧ<��x<5�!�f���c�������1Xê	��SV�4�4Բ��^{�O>���914D_�:6%��雉&��%ǯ�>�=��jQ�l��M$�����	��ǜ��p��=B�GI(�KV��*z���ǆ�ɩc��9�o��ݞ������֌����|yD�=�EL��Z'i:a�1M}KJ�?��H!׵}kl8����믻{��?d��i��{�/��C������F0֦j�����?�\�7i������5��	��Mcc���"y�H����PcA-!�{	�8�h�o�;;;�y�MN�/P2l>C�P�3�Ծ!4��b�`3�CV�)}d�'�4H��g�5�~i�1(���uZ�����>���7o�d2���j��0d�ш�(zps���(�F�J0IM!D�Q�씦ID�M�5���G��2�u�?�����-��:��o�=�I��K���ؤhQ��Ib��d�����K��%�u��Δ�*�Ϝ�]��#�9's��hރ8��
w���/>g>����a}|pz�G�9�[��B7�>���6i�fd�D�֭���K��9��6�"G5p��>����q1?f�8�i�w	P�b4X��Np��&x�:�Q��ط^g2������[�n����P-*�T�<K����a���tJ����k�k�6�k�ܣL�?Jm2|}Y��t���\��n���b���b�QT�d��z��������Y���{.�Ϙ�X��Q��s�w�i����T���*�4̐'���IڢVf��,�yU�3��u��9jr��r�����NL�80XG�ΐ��)RhI|^!HlSI!�F/��81}��;�.R8�MSr��^�Zˢ��b������7�`�X "�f��-��� �U���	wՈJ:m������A9�8g:��'��{����o~��X!�)��lE���z?���ͳt��H��g���MU'<��� �R�Mc�0M�}�6�Ir�:���rvv�x<f{k�FW��h+�8$��U��ǧ�/`<j鷼 �x��7h��DD�N�\�牠�T�Vz��*�:ùTT2������cDb�:���"����(eKW�qqq�h4b<��s��/EQ��̤ȹ�W4ՂW�~��C�����;�Ai��!���,F2��P��d9�h�+r����Oy�w����.�~��i�}��%3"��7��r� /2�s,�K��a2�є��o���8
/�P`���6�tL����<?/j/�\=�X�HUG����Yx�'�ߣJC�RH���M%Հ���!PU�шpnd.;5�90�F��;;�Z/.�*0~m��;��FM�S��1C���Q�*X�#M���d
��H(PM)L�9j"Zg�=֮1�A�s��Ⱦ;7UE}"��1@�$ǃ%D�
>�I�+O+ד�c ���4�Q�B�TƩj�e`2�$�SV&-Tc�em$%�������jj�1�&�z�'�|�/������є/;��4��}�l0}�u�M)6��o �������38=9O�![�rA"�jA^��.�����K���xe'��+�<�W����yxxLY�lo�r2��d��*l��A���/�ě�9S��bLd4cd>?#F�2��������4$gOk�@'�mLj��BĎ"�+AXGT%�@f�I�8=�9��t�<Z�8���ON��~��Dt��d��vm_�]�ܽ���ng���
���!�jko���bqq���HY���
92"��Ĉ+�;W~1s.o#Sk��r��}�D�w���b�QgBPT=���Gf���.� ��D�uf�1��)��TbhpbPIE ��!�>`2�8/��i�e��%��;�� �Tu@LҀ�@M�l�bO�>�+Fi�M�eY�R��c���8�O?������K/���8��g�/{��ED���{��#�n2�F����9��޽����z;�!yF5_B,g	U[l�f�����_����ې�T�"�	��TeHT%���t6�Xt����o*���y/׷=!�L���,K���HӔ�u�d��e���5����]mhؘ�����i�4��jA�@̦����]f-��kV��#՞�vm/�׷]U�1\�e�p;ϳ͞@�Y�X��1�A�TU}����ON��?{f�/�(6�m�bl#"�����L381D�k��✏>|���}k_.�W+��QbML��;�o�R�C̞�Da���e]�Tu/�m3�3��&���j��0T�Gu]3�����{���9���a��������g6���#b���]�}����\RUu]����O���S �˫�rw��� �qA�\�4�@�T,.��O�WDٮrD�d���>�z/�ʲl�w-���ޝq4>0�888�9��E*�0�~�~�!����[=�v}K��H����ΰZ����g���G��%w�~Ip��k��9::i��5M��*�
`�!�P.�|�f���<MN����d�x<���L�I]c��c$gwwc`U^�喦IrV1�)�l�Ř��X�\�ָ�F�awk�r� ����M���9a���).˒�bѷW792�	�k{{\�4�޽��⣿zO�>����yHS�g0VԊ1��)��{��w����z�c���=��W�FFmQ\�DH���N[�,I���L�,��pbhV�|�q���C>��"7�/K���'ڔ�M�����(�jY��S#X$Eq�U]᫚&�ӗK�UU���!�oW&�e�{��a4����*w��q�rY����o��EU���X$|�J�z��p���e�"�-ւ(�� !��^7�>ǫk�?�u�W�Ɠe������ۯR�%���#��Ƭ�ˏ��w�e~r��"bD��Lr�o�U��y�l��Eç��\R�O(�r~|ȯ�����X2�pn�b�"G��ܥs���4	g��"�o�m�c�t�у�Dk��L�,U]�\�S�Y�D�Xk�&G5j��E#B���qD�4U���A#�g��k)�N��f�v����k�8��ʲ�����qxm��U�c_�{gO�?o����~�b0F�5��&���n޼��ō�)ҟ�=��w�������)�-�<ʺl��1�5�%���5�bI��3?t<�x�o�ۭ"6��ǋG�9,��W���8ɋ�X��M]VU�Dz��\8�E�C�V+���\<M㙟�T��P55�npy�"�F�bZL`*� z�K��*��>Pi�f�RU�,�X��e�ȋ0��y,��Y�q)�g���dY�V�n��B�W�$����6�Ʉ���s��O9?����b�%��CįR��u�Z��zYQ5�De�8C%#����/>~���C��h��̦	b@µE-�l����}� ���Quiq�7�|�;�����cV�c���L��V%e�b<)���Q�d2�ڌ�+U��TR�dY�u�H$���
2��Z�=�1_��>p��.?��_��_������Š�9L�1�u�x5��ڮ�쉩�+
q������:&�K�cH�"W�5���S��oϞ�X��k��Z� �HTU���|�ѝL=b��G������:$3HV��Ħ�g0i��M�n��ih�y��o���%b��X���w sC���W`\DB�$s��ƈ� ���Ȃ4�4�@R�h5�h CTPb*&�*�T�8 �4uE��T�+`MFf�����p�����E#6kٸ��9HQ�<Ot:�ł�GGܿ���!�Zsc�(�E4]G�,����t9��H�o"M���fd.c����(9;:dw��l�x��t:�Ν׸��Ërp�6qB�b�6#����c���x�s�h�Ay��7�ۿ��|��'���s��U���kϲ\`,WgL�c�[3D�ղ�,=1���8'+F[$�-�Q^P�9���9��;����bvp��;�����Ǘ_|�~�#�#�f�Nߵ��ܷu�$L��w���'ڷ�1K�y#��c��2��o�[�N�ט�?{f��v�:�b���*�X��7:��|Sш¦�}І�dy�Ү��Z��XMU�Q#<j�t)�0Kǟe�d:����m��2w�0߾j[�+-�#�Z+�#��k��P<!`l�o�<y�J��u���I)
�!�DJ�V5�¤pX��@]�I�t�\���U�ˮ|�Ҹ]�9�}�z���)���dY���>�W4�N��P����9�t�Sa+w�Y>�19���h��d�l6�ƍ�e���)[�F������wU%�e����.Oc�Bh��=Ս1���͛7����;�&PW��Δ�����7g<.�
G��M)�-��	�%�fx��N��bB�;l+?hPʺag�s�/jƣ���h��rō��kQ�k�f쫜��c_Okݤ�Z����c�ƈ���Bhv�>���GnϮ��\�&�Fk��Թli�� ��4*D�Z��0��n
n�U��S 27�p��h9PhkNr�VI��AD%(fc�G{,�����X�i�@;�]a����nL��v��k�1�y5o�,����t��
:'�;��HL�A#�2�A".��?��Zub]�2�D��q3�����	�⮃��n;��x]{w�Q�z d�fL�H0�&V�|L'�r��9��.+�嗼�ڏ���f[�ᢺ��k�1�@�R��&E�@�b��''�l���MB��������bl8�4~������t:��{wy��O�h*��7�M�Z�@�'9����>� d�\��_-ɳ1�2�8�|�v~l��y�f#���!8�h*"ڻ���N"���=`���c2��뺯�"�7����2��Z|��0����ވ�Ez��L�#���YY�U8kɍ�=���>��|�/��ⵢ��:,[z�W��1�JQ3������ʠ�x4cȓhyb.,�^�~{�=ɋn�	��(O�����/ُ# �t����ߴO�� R�} 3Bp���E`���Q��&XS�e��UxW����?�y�{��5��OĞ���{S䙫�1*>Zc��[b#q-���UX�a�eh�^v������.��[*i�H���ገQ0���V�&��ld�1;Ƣ^9�H��!�n;,���E����988`6�Q�k��,���L��~�mn޼�;�ï�ׯ���ҴE�`ggg�6�,�ma�e4�A"�/IIB1��\I<b4U���k�:M�}�1B�5>4L�#|�F��������`2���$��U��Q�o,1
D�c�T�h�(��`\�ƫFa2%�ؤIAfZ̆���hDY�,�ˁ��z���i��4Mr>��#�Yv������o2��uXG9�e9�*B����},Յp���gv��E���K2.�2hC ?j	��ݴaz���u��/�Jr��].�����I�52t\$����!JE�%�����?g�H���h���Ísꎣi�6ř����-N�N��S7%M�B`kkь�?��w�}����_n�\��'PV�1�,3��cb�+���Bւ���K��ڳ�͋("�!�,��|�޻�f3�g�̶o0��߿��=��%U��E�t��6�x����o/��yJKR뀸Q�~z��,k�j���Q�1��.)˚����_��8=;&9Ǯ'��a���x��]!O*���Zi���x�i �<C�Xk]�qbȂr�!F~�_�������OĞ��3��7�I"�1���E�T��=�${����m�B�N�l�L�pi/n���f}�YqI���rT"Q"Q�zNY/�}�ƒ��SV��ƹ���h��|� �EU�V�jA�G�N�Y.�NJ�+֦������"b�1pcg�<��f�X���i<(�3v�ʀ�a4v���INP�K|(���
Vobrh�}/��M���O@TT�s_���rt|�'}���vw�x��g��z$ɲ;��9�^[|��-2kk6YlvOw�C�%B"��a ��[�#�A����y P�<$j��iABJ�fi�Iq��j��fuwUu-��ofv�=Gf����UDdFd�/��%=�����=�,���ob����loo��u��޽��l����x�Z�qU�ށ\��h�����֢1fޖ��*E�r���>{��t�<O��!�������-�d]:��xɕ�=ǵN"�u�:bb��u<�����t��2�܎Sd��I �@4��j�U=��dǵg�*��tQ�Fg��f�?�"@Ϟ=�t6�phaB>L�� ���SXAVa���H]U� �AQL��_$�'*��s1���Q�ʢ�?Z� I-zY��J�O�0@N�1B�D�"v�	���w�q����CiP-k� h�	�z�]0��5��@9�FS(����� "`w�)>��
U��ܹ���h4�[�-�R�4�p8��=�y���~}~��ԲIm;�v��j���i�����柟eOD�    IDATB���rV���^
k�n����BT�bTUk�s�5�P
���lx��A���Y������ z  2��Pa,�)�O��	x$����&��d콟W#��*w�2����X�9P�
Fl��	9!����e	@��C�Z�n�����F;�L�_�V����PI��=,�1�e)����
�H8���3T3f��k*(��H���D���~��;����7�	�����!�=|���;��U�髯��誥����4 M�
�bŬB�B1��5��0������a�;��$�F�3uol� !�ab	A�6�k�I�=��pi��u��Z�� e$V�������1�.��s�6��x��9��)� ��|�s���e�䝄��'Q
@��a��"�"�,S��͛W��v���W�z/!8%�* D���(����m��������
ۖ�*�8Lq��w���һqR#Ԇ>�b�<ϑe(|T�߸��~�����;��t4; ��\=<�H���$I��iӓ�����|.�=�L��o�7n��H����^�\�=�=���;�ֻ����|@ݲ�52$��X�D�u�PS�x�������b�B|�?�s����B����y�$"F�H���3(	�� �`!^�� �����E�S���ܓjc��U����	Q��!��7� �Z���Q�T�^�7n��t:�{�F��"��hpG�kD+aԎqQ���2�<��n���d���~`�k�錾�z�*U��V�B�D�(s��{�XΫ[�������úz��W�p+颵D��AF��`r�JE�;�o�w����.b9Äj#�(j� I�y�d�=vvv�OZ��s�!�j	�,���E== �L&��X[[C�� �3��>���.{I�!1)����d
�dpFPU� ��B����AljA�3���*�:��	����g���� ��>G����p�]�k�
H��
��U���A~��c ���4��i{~�6��Dh�Pfn:�� � iB���I[lT5������1F|��g��f�y�fc����u��\�H�q�ڕ�"9Q�(��T�bϕ�1��_��\9���'�1�5�� �����g�U�HI�`�=�u�I3�:|���"�<:�+�$I%Yr���4�줉ʫ
-΃�>ŋ��X��D �ß�uv�"���XW�Ɗp�7���W��7�o�c�����7Z�+�v���4=�Z��m�/�~��q�1l�s�w}�[JD��p�U�M���d2�͛�P`2.����|���
����A�A]#r�Ź�q���n��|���`!�����)�ky�Eч6�#Me1ڟtt!w� � �}����X��펡	o��%�(s�&4���RK�4�i�@u��$I���������N��أy��a���뻼�Yu}~.ڨ���q��w�ߟ5�q�y��H<��,?�X�Ԍ��M V�9��9�z=$���g���!�4�T�4}eP\]���������������w��>@������.�{�ۿO��v��kU���p,�u$t]����q��[���)qD����S3�xv0b�x|S��vt�\�
!>/.�-b��x���,��v�B��ԤU�DX��a�����h�V���b|_Ǹ����o��Eh`�~�Wu��A��w�Qp�kG,���i,����݊Dn������PE28*A����=�TM;2s���|Z�r�Q����K
��*n�婳[e4.m�1�)���&|׺H�̊[[�uo��s,���풂��L���cgf�S��f�Zs���O?@٦��n�´��@���wtA�3?����i0�3�f1��)�L����N�
��x.61�� �C��$�a�۽`�K�Y!����D�Y��8�p�Ԫ�@�>t��Պ4��Zԅ��5�.Q�������;�����q�V⊄��ەK��g�R�4��o~� mf�ciߗ�3��`8�������sW����g�$�~y.$�Dishq#�ڻZz�P6����?��iM^'��>U�)�������VK�>����Ͼs�G銼�d�+y���n|J�k���|<fn% �"������ ��
�K|���WB�q(����"Y��e-�hM��Sm5w��@1w�&���%�>�q(N�_,�ڗs���^m�_�1d��F�Y� hjd̞E6F�����E�<�K���R�İT����eK?�t�*�r���)��w�X�m�&B�d�5#2}����ü/�m�ZZ)�>���35�_�֮�9����Oj�2'K�Y1	ͨ���Y����c����u����U۽�jl��܁��|'\C�UDJ���DpD(b�/���[�����q ~�HJ�_�I�6H&jjf�p�dBI-S�q��*�l�H8�����ڍL��H#p���o�OX^M�x��4V4�_'*tvWI�"�Y-hXT��"���?�&�]w�ͿMb���չ�+�C� � ���۝&�m62Q��wd|g�����Z�jL��͛�$�q���J9�eV�����d��{*a�bЁ�O�e����l�2{�bu��2�P;�z�݌a����ݿ���q�m�SH��� �n�C[���f�F�Jg���h4���*�𱱣�Ш�H��	��U�;A�0�c��W�B�������MqX�մ��!���D?*m�0�`�`YMa$E��g=� ���9:���W-�%��%�����1����6�+��L�W�%jf/Vu�0�u���s*��
��
�w5�F���v�e=����{Y�수��,�5*a_�j����*�j*lU[��P+,س鴪�9��y�?^��p�Z��>f �E\�r�"��Xq(�Z�k��}e>��Bɮ�V:�k���T�"E���8M%�M:E�i�􅲯B�ǰ�*=�Z��O���Hl8"��� \V��:%.y�����t�Z��_�g���V>/��W'��9�C�����Sc:�.��O�_��������ާ�9�ִO�_ZiѸ�	!ı�h��_��\�?���Y��I��W��G��}�e�h���[�������b�lQ��o����R&���E���Y��u��;�#/F4O&�7J|LݽD�:��\U3*]f����0�*�W���P��*���}��{ c�X%|��P n��1T�W����k{��֓��|�?*�{�Z[lO��k{�׿1�g�%��
�+Z�_,�Ԥ�Z� ���^I)k��g��(y:kƭ�N�ؠ�O]�j��j��HK�GөzGǗ�������B�X90����܁w���`{i&a,+;f>j�h����d'��%W�Qk��9�L�W�' Ai�gq�F� ͧ%�����f�u�o9.��)A�ny�_��<l��w(Y��4}A�^���h��ύ�6�"��`.��~یl�Kk�D:ퟤ���5q��l�e�:pF�� i;.�A��/�3�SEu�*5�^���5cC��~dO�^��S��#����֒$"�*�qP�7�o������yW���WM?��o�rMcu>�tJ��.-����x>dp��|���?�Ό�z�fَ��9p�+�̓��DPή=mO�����\�7	�FF��M�Ց�Tf{��RKE��:Z����<{k�����o�{{�B{.���vߞqU	�in�P190!΢miL-�O9j�a7h����1�}��z&L1�IF�)V�#�)����!��4v�Y�Wn�P#��P���%���.(���VCϕ�J6�=�T�%d�*�+�f����e�=k��Kj��צ.�92�6����
���a9�d����Cz2.�@^�QoP����)P�<+'��xE�'��=Md�;.K�E���x���l�HEt��p�!��O34"�:΀7M�sqlD������y���d�XN+�I��%�u�<�qve$q�RRi�/��4�ģ�o��XkF	�E56R`Vh�+d�K�-�t�s�S�6���mK������jE<r˳���C�,���\��P�Ilf�;�. ��g�zo,�eTE3"7��Q�Zьm��n�����P!P���a׶��G��3�B&��rK\������}�������GF#�����{\��V�D�Zp�/+m_E�[X���Xִd>��,��8呹	��l�K95�~���ңV��sqC-�H��fh�~����C��r-�����̕H.js6��S>[;��"�(hmB��%<�M��u���+D>����
�=�Ѐ�˱���,�����0� �o��D�	X���}+�$IIIk8�SW>0{X�%����_���˷M[ �}��S9�&S�I�������9�����sN���|��*!�4b�a���L=_9^��$��ys��q��b/( ^�և�>��d;�����d�E�T{V��Q=�r:��l"�Ft[Ă������9��Tg��/�����'����!�Yt����!�YMG2����p�´[���QDJ�AM|J^�1o�}�ƃ| 1'�!�7��G�7|/�X�C$L/��j?F~��ώ�'�IY�gã�R�"�d�d�ꆠ�:Z�ĝL��?�}zS�ëq� X���λ�VZ>-�g��Op}�S<��	Ƚ��611�LB-�K��v7}��탿��1�qq#�۝��]��*y�rF1Dg̽%�ʲ|�Tj�@����z�\
�~z��66$@Ʊ�DՒG�_(SB�d\�`2c�.0�=|f߳����W�^�j��[L��#g�"���t+�X0���˚� A��3u��L���|�j����C!�&�t�D>,�Z�t�������)��I=��C@��ǥ;��5�}:�}�[�h��B�.2�.�AR�y�!n�.��.\�X!=g2�8+�ThO�Rj�:�¢1k(0<���B���E�H��2�!-%BχŀZ�S�h�W�>�Y9��_���$�i��o,�=L�y�Il� m��8d=F@'�|HR�`	9��P��{��8�srѥd��t���\�ċ�� ~X��ݝ�3˔0�-�͘/�J��O����x��ƴ]��[_��G���v�t!lUP�I�2�u�/D Ք���L��(E�LG�7����bZ�\���ȴW5�,�\[pر����qد.���y��O���f?l�o=�~E���}�F�����>)�uS�e�>�����sڨ:TH�_��m����E�$:i�]~Ft�zҸ��p6a�I���Z���:u_��,����h	�A~sbR�U���~9o��E�uN�g�������&��d$R�4E+�9R���Xȇ$�/��W[�^wMY ���DY��aG�}~�����}̓�>Қ��o�tn��'6�.��`q@��4�@t����<��J�f�rMو�����1 e����Y|���z��{7�옾�Z�o�����:G~jK�6����TM���f������f�LF@�D&lX�j�1�3��Q��NJc��+1
�EL(�Xj�4���_l��C2H�-v.�������x(6���N� CJ� �\0�Y~j*����v��`�n�����3NRlWR-����������T������Ժ���WeP�DH����$۵��K7]�h���9�5۠�܊�����i��[/��.?�S�0���j�~a�FY�	<�Y�kGƠ�?��+5��@|��`�ge��`,VN9�3���$O����_�����q�Q��0I��Y�_&R'��K�>zF�
Y�T��i`G=�ĥ\�`����~�x�Yd��i]e��� vB*5�$;ﻩ����\��$\a\�� ��4g�Rj�V��\#�%%�@��|�P#)��q������8�W-����q�p$,�"����%�$�/�#w�Q�!���>���G���ĕ�C�~��'� ��޴#�&p� �zg���S#\e���!
��s:۱Hi���DT2R�������0��1���0d���ԋ5|e�2tvn����������������d����L��Z��2��1nf��CK�hp�f	;$�K��^�W�9VQ�1��r�u3�u�;��S��(&��	je��A��/_��Ӗ�Ц;�eP��U�[��b�A�d���1�����5	<��g-ԕ ����_�x�&���&hu�чe��]Ģ�?즽w��:�����]!� ��7�֎g��wGPe�M�����8��׬>��f�P��G��(����Z��k0�_��Lw�����'��w������ܸ
�gh��sUceLM�f�M�5G�g��ݙ3=�!���Rm��v�K�׿V���%~0�VPQ������P1��f^�,��� $hf����,{MkۂA�?B�y�X5�9׆�T^��}���SAy!c��Ie�������,��K'�6LY��2�z�+��Eمϟ��Ѿ��<	Q�����A8�1'�+��j{h������2��K���C_�(:o����������=,~���X�o�/i��~��ۧ��sW�a�`�@��M�qF�u'+)郎J��	��n�;l�Q������7��P{�:�H�-�Le�]���?����zo���@#����x����X���GM�4+����99��PX3O]���P|�Z
V&�n�e��Hӵ������.�ҡ�`E0+�i��0�}hq�.�
������0�L���n���/󾦫Kv��]��;���c���ZON����ޘ�������)�Sa�S������O��8s����_��/��������D&��v�[��v��{���|e!HN�vWx��3�P�lwq}�v5��V�N���-�T1����7�w���SߚF��{[%�̰x'B,^�G���N��UZ �����A��q���^��
�)�Y�6���Ͻ� [�������zݰ��	t0�QP$�W�l�lu�W������f(�)�Oo,>E�!I�����!��g�bH=2+ǚ׳�Jg���sC�e��0�)G��2����� ��6K�ڭ�P��;���@�2��%���p���~9��?tn7�Z����m4q��ˇi�\F���PzׯT|�\�J����K ���p^�H��͕����t��Yā>�qk��d�K��&SX���Я5����
��x>ێN���3�!
�Iy��oA�M>A!���:_L�w��}��8���H'�
r��=T��U��B9#)o���:��'>�;�)������z��Ҥ��!ɆA;K�WT~V� �VӀ��u奔T�[PwY\���ڏ73���A8,������i�!>?��r����n��g��̼Y�� ���qbuZ%���4�){�?T�@gQ�4|¿ո��`���c[V��4���i�s�������o��/�,�WN3��C���F8#(�l)�*��U��_u�5nZ��o�c�Du�&�[�z��O�/���}ă�ݏ�}y�>�?����u.ՕR,�1���N��Mν� .n�SqG���d�(�M�$����#^���<<A���͇��n��M������$�����x),����"L$�V�g���&�Uj�؋@N�U����������܌H�s�/����\�E�����moΞ�˓��:xm�WG�83���Y|�H����;M�:JU��r3Ҙ&�@$��Ÿ�y�a����2�:�4����%Ȓ-� ����tb�00��
�+��!�ib@���{i����ܬ�,H͇�j;XM���I5�?����@�tq0�U��Nx��i䕿g;'f������;�&/�֫Yx��DG5�t�I�p�;������e��"l�}�]�b|[O*|2��&׬Xo�"d�H-�����o[\YBv�|�o�7,�(�sh#2�T~�ڎ���3Ko��,�IH	cr�C=\n̩h4����Dگ�x�����-�'�"���k_�ٽ���"S�k�zW�6��ab۵����fK.�I-o���X7�)ŷ����U�-��Z>�v�|M7Fh(�U��tj\ﳒA!be�APt{�/~x��Av���=�^�X���XL,DG�'���G6�8q-�̧����@�m�0y�^K��������EG�uM�~����w�3a%�������ƛ������LO�g��n���n@*'�Sv�V�I8�]���.&NǞ���ã"��/��ؐQ$$k��s���c/���(x��J�յ�Ⱋz3l�G�RO�j�Wb�(�#��X���%A����o�&��s�b�>Z/�.�h�_��W�g�Gy哒!a0�R����7�g ���� �0�@�,�n�"tg���������)�+��5r<T#��ߔXɵ)0?Bo�F^�-�`0<�@�a1b���ƣ���i�D�#>g�1-�膷��j���.$�-4�����}�Á��{��Y��N���[kC9�퓓�	gj��FZztZ쌼���2����G��̗���\l_ϣ�߷��'d���Dh��m��0M��T}�5�#J*i�J�w��Yp�%����k�5��9^\�O��U�rt����rKK޹�Pm���&<�(v��+t�2<cJ�Oƴ}���9fg������4��j���ʚu$nG�
��џ�O���u�aJ��
��v+�O�GQ�����TVU-H��)d��֤��*�n���̳k�*�T�Z���.�5�x#E�4�c���L���I�|�*�/[H���C��G���^�*H�'ͻ���U�)LC��iz�q1C��o=�e�o�}2y|�3=�M��U�QT�����ݲ�L7��\M=�zmXw�c�I;Vj�P^4��e�3�S��/�Ic��`:���_���h�~sq������u�ϲ3/����v�<�?�NED�+?Zߌ�s �N+D�I��(�wPD��-+�$|	Y�g�$6+��.?�Z����t�3`��<h�Fru�E�K�qÚK{w鞭v��
xF�v	���"���P�D��pJ�Е鉜i�r��g��&��Ʌ������pe����'�w1�A�X�JAV8 ��4̬�����O5��_�89�?P���w�c(��f*�3��^I^���L�{M���
ΜO����n��oϪ�c��^��Om�?[we�v�6�������3r�w�\���l�}F����z��׿��_6,�����oq��-N�O��	���&j�S�\�Q��N[��X�j�xवc�<|���UИg���]=Y�s��`Bx�56���l;n��κ\�9��d}�/�'8 z��MNO����k���$B��u�qiC@��%����1)�F�~M���A�����@�����`z_Cn;]�wI·��?I�`\7�������E����d��gK�����1;TnG��r<���J���H��Ժ���y׽��j{�H��(Cfd���o�K���;^��9M�@�CS�����>�~n�q�����S蔒2&V���1���^�e�H׍rĵ`^����M��1�������z��E@Δ�-/0c��d�P�7EM�����w\\�h���&�����g�@{�ȧ�5�}����:��4��Sf����f�.�+�(�X~�/	��_�Ǆ��lJ'Q�4��18±<��+�_���	��<H���qo#����?MŃ۟!��7G�ɟn����ݽu��	"��m�cO���[�!/|�����6�;�
������y-��T�v���z7�ĳ�;��G��CPx(`�*!��yY~e>B��	��l�����{�H�@Ҽm���r�'n>�;nő����0"�F,��@��򗑨�Xh����Q�T�kZ�f�Q�Ol�����I@ȃھ���$�{� Ʒb�n�M;;��@���xOk�3����z ��o:��u�a�O��1��d�1gk��v�J���|���2�  hen��86�sJ}"\[.�+sL���}]�T���$J�+�3\:S����{�*�	z"�8�|fA�2K��.��긶����ո�3�M��5�e�x�|OƝ$K9Q���.J���F�6��6®0�>�
�؏ �{Q����q�oh���!M��2�'y��t ��V���Zy������򢍛����Vv��L�� �{.�3�7��� g�1y|��|g+W
7��	���xh*�s��0���T�w}� (rm��ӏ�b��")��k����JT��p	�H�����8 S�9Z'��B� �j>�DCN��J�#Lp�HlS�$*�D�'i�� ���#q	�$��W��G�ogfE��w�t=���yI���dbb�DS�c��9g�˰��n9޷c%����fb�(�w��\9����n؛��s��zF(LV�.}r���^��^�n{��vݴTX��jB��P�gee�e�@My�m;�ω���)��xy %�������)}�JO��?e�`ᡰz�,�D�VZU���o�Nd~e7��F�V��	�./j��ܲw�W�դ�����񅄈k|�*bb�+\T?�˟@E)�\y��h1�EB��'ؾ|Y{ۓ A���Ɠ���wϽ2�F{����aƶ��iɘtm�E���s_�&�_�A5/[������o�h��hp��ϹJ\S���7�";���ʡ�ӝL����ʙT�����L6R�I��r���l�?bA[̘gY�
Y�7@=s�P��Dl��ׇZ��W���K��!�=2�&1��G��6����h(�?��\�c+��R*9��)#�H YU��y���>��E_;���  ��f�j�e���Yョ�ޡt�x�_=|�r�b�
�7���T|'����G�
8�E�,^-��\����
.n�ӷ�5�A���z_!zSO�宩�f�I'":��������H*S� 0E���?�}��E��_?�U���7�W/�Vqf,b��L�4є`	M"�/,|n��	�/**��f�ṷ}w=��,�+fS����ᗛ���K1��"B	�ݎ��5Yw0��L'����:���k���`ᯮ6�4�W�s��X^��Nط�ѥ�^T��vPSp�<� ��iU%�����g�MFu��4��]cg�-���iZ`�K�B8h��`�����u�&CJ��a�q���x���b�q�$�F��]QE���F�A��T�́��2��F��F{��i��l���/}�H�&x�@+0i���s5(�us2?3r��@F�B(G�o�=Ώ��E*��'���Q��SǷ	�����Z(�X#�"6����y����S�IE~J*ݤk�O�t&0w.��O���(ͱ��0��6W.�A>�����J&��lM�6[v\\_{up��F&�A��@��ꭞ�,#�M�� �W���e������c���Ǥ���3�H��j��Bz���NҬ��v߾g?�:�N�l�W�U.���jp�59���
QMѶ��*�%��x�cn�u���"j�<L���гhtY�w*��$*�B�Ԑ�RiԬ�(x���hh(���vu��͏���rۀ�|��_���%�<V�JI�L��7_|O6s����mЗ��;1L���������㿖�{t�>�,5��?D	�{��Y�E����RM��� 5 ��܍�E&��M���UC�!j���d_z�_����ƣ��`d/�\ݭ�_7�v�q*���Yt��C=ӌ~w<Ɵa٣5��5!3�Dj�A�J⧃͢�5��8ס���yՓ�X�$$Tl��#"��r
�?v��5=�c��0� 0��!�"�ՖI���í��)FS�&#��CC���YR�r��-������H�\!�r�9�+|W;���h�2�j�^���ү�̨55S3��x2!�y>f�B�~�@�A2�,���0"�h��	�����IB��@Q�v]�rGH5��eZ٤�5�����\�����E[���2�j�|�A�k�R˰k��0u�3�A*�r��}����+�߁���3m�-���_�OW6t�����7lR\6�gw
b�q2�tJn�]*�X�G��;��=<R��~:;s��q��D@�8h_��10��1��y�Vl��.Q^ۖ/���uo��s��מ��T	��xV53c��)x�e�W�V��A�� �j;�[�h�7�(xo����5LEVk;��u�}�����<���HI�
�Ї�^�@xq�C��d��8/K��*q��=L�pkqk��g��g�Bo�C�k�B���Y���G�����/3D�\��v��}�cTs�"�my52�M�@�T����Ǽ�܁-�ʋdݐ����=2��v	?x��g%�ӯ�_�\�5��#��gU�j)�ȋA(�yS�g�l* !_�]H� �i��S�qs�,��Od������e-�;cFY����'�2�j�޾w�x���7��\騿��ԁ���V?�.n\�s�Z	MJ������5�I����>8��B���w����7��IOg�O�pG+���A��J�U�I����`*!��'�G��Y�p�0[�[G�*˅�}������4���1���N{����
_�Q�q�`�V����"U`*��g���wm�����o<�nٱ/in�&{���_P���&�Ʈ��P"��bg��(xڔ�B\FU�s�m~�����n���I�'��n��|��#U�<�>��T�-K�3��Д������SB
��<����2-����Z.���0cY�hZ��7�m[���X�K����͐�iu��铍$~Ԥ�Q���衆�M�S	(Dܾ^޶6�0U�^%�����'���n�=�0=N�l��T��\L���$l�����bM^<��ʥ_�#@!��&�(���8[�ވ;��PV:�1}�Ye"��K.�Sx�8=��
�<��tC���4��İ�j�$�B�|��	}u,A�����O��mc�B�T]��;s��$8(e��Z��j?d�q��6ӌp�#��\1?`l�^#��yÅd��Q�ح��Q��R)�g<M�@�ϵ(y�����s7�N&�q-jY�~e*�,@!
�*"$�I!�/�z5D9���f�ņ�l�Ww���68jڝ��0�K����*�Y5�O㨕*{�� -<�&��dX�^fs�:�Q�����_��&Fe�fğ�J��ۺ�I+�rp�^�܉�s=e;G�����`.�
w����J��q͵:t,l�P9�>-ڄ��	����7y�o"L�j[:���ow�s�\������HR����K�#&�K`N![^�C��LȘ��,؀v�%2$7>U5�������d��gP����Uu�6aF��J^� u18�����^�uTDxX�b�/�U}y(� ��uh�.��if��J��1P�T	��CG�ۤ�����*���M�%�Df10��E�����l��d#���5�������
c{�<5zW	����Z۝�iB�#�X�H���	--���|�����a���0o{�$SYm�kk��Jo�%�����
��Ad1�d'�{ƿ��g�L�����}�@���	 ����P\��pȎ�k�Nmuz�|��N���wnd�l�5��-���D0�%�L �T$�J
1F�%�����&���mGx �ƚ�հ*TJ��a��%?��SW	��檜�Y���3�!=�^�_����9�Ʀ�R/ɊO�vU�v��Y���K�߰Ʊ����E?iW����֠�%S�%P��Qa2����#a���#��uA����_���[�{{�Y���I�Gc�0p��۵�KX�嘼1�j����M�n��rYrl�����C�� iZ�*�o"��s3Ɯ����C]�������Y.�����=~��������h��h}���P���r���&>B���D�A�?ov=� &r
�o�!=(s|�g���,���ɀ)��A�jր���xr�Kޗr�!����~�u2�-˘�����y��g��66S�>jq���SaIY� (��:%m۪ʔJR�G9�X$b�ԩ~�K�Z`���[*<���W�D�-j
���^vĆ�!��>o�Jph�Ḛ`@��,H}��@�?��9E@'����g�+���HMU�.�)�5c����hC�<:ں�b߽i"��q��3\�h�����{��Ǖ���#�� \�~ؐ��U���zv�V��~�A�{�_w��NrM��&C~gn�C+Q���b�)[1�HD�G�G�΂���0���c{[ۢ��m�X��Ȏ҅��bP �Hi�Sy
�;9��"�W~�	S�
���m������A+j����sL��}\��D������{k5 yxx�&�?��o0���ݧsl�X��
���&Ao� �Y����7���:���,��M:*���פ�Gs��GA~f�Fm�1^'�42��yq����d��Θ k����5������[��,資�&FfZ[�=]Y�X�*�=#�r]�5pM����-�y�嘟�������w[���ލ?Å�I�>��(�hJi���3�+EjU�ɨ���'J��%uѦ��Z空�����n���eu/-{�դ#�5q���7��w�/,.fD3�`P(E@�����ݽ���3��_מ��k?;1���VW�2�ĕI~�p�2EAO�~2	od�?���'��N�+��܆r2�48 �~� A�%H��1��1�L��T�֗a4q��~�r�v|�o��4!T�tU��GP˛1_�؞ߞ�w3U���ԣ穀<Ec�"��/	���P���al�T4E�����ݴ���ܘ�5�1Y��+!z�:���ɋ&:/42)�����V��3�t�Tj�*.O�F�\M��À��*���L��K�*�w&�	�[l��H�����7���W(�B��?ц����X�w+�y��#�)O���GQ�>MSCq|��GI����M���뭨;)Щc�E�	��j��[7�Vo����	��ʯ�{w���b�C,�l��E�����@�3��j�-X�~��_����!��r���3Wq:�wI��7���Ns�|I��^�}�dO����$8�r��v�̊�H���p�c��7��O�+,��Z�;����y�7LN$�K*��IHF5��|�@<?�O@�8��o�g��z f�6
�����'.���/S�Ô�l����<���;ã2����,£Eb1f�V`��T����7�)�7�2vL���+��ŏ �������xu��@���w.�`F��<�$�#�h�:U�&����M O��T�Ğ=#�̫H�LE1SI�k_���}>���H���=�g݇�u:�ɔ�
���}���,���w����B�ϻP�I�*d�y�\qX�^���to�q3�a��`{�%���z}���sWmt C4T�OT50=LR��-�\Ǐ����ͩG�?�#�J�ɦZ5A0�t��F������y4)`p��*Ԅ��{?]Yˬ���W���ge�T{�uv��g����t9����˄�5:�A�^�=�(t��beK�4�l����u�6�j�ءL@������eU*S���vX����d����OjS�S3�L�0�:O��"��=w/9���~6�CJ˭�Ic��o�`z��{ϡ�M���g�vE9���wX�1�M�!̮Pm^ٞ����L&��"c�"�t]B�j%{h�����Y"qlG�@"���o���e�Q�b%!!!FM��D/�)�9���(=�/p���+ ���ږX 4`�?�����e�g�\�i��+S�k�u����;�`�.��Awl�D�`|L�Щ5�
طBƙ;G�׾g��G�c
x7?@.�Ն�~���h:����KjKYI�/	ɠ�H��H��S�҉��d��Mj��9��
��v�Cw�JQj��w-?�ne�=U�3T��nF�	>	���@q�M�b�*�_��<GlO��>����R��iQ�6���?�N�|_����9��顦 ����R�*(�f@���Qڿ��6�έpc��D�:L|�o�P�6�|�{-�y#;��Mi�3Noyx������k�8���$��ּꜯ�w���k���B	1�#Bm	��qp�t`�e�P1d��v�P��5��	�٧z��Y�)X*��bD�|5�����3��gS����j�Xb�z29���Z����"A�����7^!��M-J���1u���4q7����&&vo��W���~,&1߇ q�u�l���ۗ'-�]_�RF���Y����H������{	��3���]�yp��lk��g�3��$�[O���OJ�w���k��x&3��q�H�,At �`�a!Fb�[J���z��ũ	|:@4G��9�OR��0΀��Ҥe,&�8s��C��^��;��@ׇ�,���D��I��@=�Yo�q�۽��ΐ��`(�sG�{��նVϗhv#u��6�.�S����sU��^��X�}�!�I�O�Ԕb$� e��YKz?�̭E�c��?妥�E"6�� @��s��%=
����#p.�� �X��ئ��\P�aE �!����]���;�i5�m�e*�������Hi�P����b�3؟iV#�ts'��7�UظѮB6��lK�����y�M҉��j�Po�������������g�r:��f��8H�H�C)5]�����z\Cߦ��*/TvD�H�V	� ���&o�������?�Q$n�5�Q0��땢�
W�o�99�[7&��`������M_�
wy]#i��}2����v��PZ�b/^�ݙt�����yt�`$��*sS8���z|��I1Q2Z��Z�VG �y����vX,#R���fX �B�ŤX�X�?�	���x�:���N������p㕈HA	��iw�d��t�
���u����_�\4�������^�	?�
�M�e�~�₎�a�ο�	��r#���?��x���x{{k%����:WDi�\����_E���5S�U�YI���/��7�L?F�8x�7t��id�Kf��]X�{�W�|#�w��Տ���B�աINT��ֳ�}�22!�Lma���~x��7�]>O|.�S�`��7_�?�?�5�z523���7VG���]dޅg����$��c���5��p�Q� ����C�a��~�i%h"���u՘�-f�z}���i� �����N�;�z�r�Է�pD� t<�8���XI��:��)��P'�	
#��F��J.�<n�FO�LN��bݢL��A�̿ ����G�Z�,U�����	�G�w��$�"�EO�C7��{3@�ۄ=%y��&��lۗ*����؎�%��]S��+c`�N�hy/�Q�?���mCٗ�)�C�&q_{�����[l��з���J)�H�d�ym�ˊ�(�
��\�&����N�)p��z_��V��~r��	�}���b4x����'J��I)�)���O#��$�\��=�m�����������m޶2I|��eϸ����gmfo��=nt��Ob��8���9�7����B�P�E�O�o���ϲ�<�ʬxQ�����g����ދ��;�������BM�kG��6�ӛ.tY~��y��}z(W1��5L^[Ȓ.��]�K����u����=v�(��p��uͻ���P�t1�ZE�!������/Q�iR��L"AwGKwC�������^�����ۛPe���M��`#�H�fW�
i%�P�����@e���3�W��t<�c�ˠ�0++X�y�����6��!�Gw�|� �J��A$a���>�v��d� ��#,,JQp��^pW Ĭ�)�����POu�Q�(w�pbޮ�ПL&�Z�(�&�����x�I@�Q���/�#c2�r?+����%A�rF�R����w�?�Tg�r_�������{���=�_a�V��������o�`��~|���p�����0�CK
,�����훷?e�*�K�Xʝ��.��E��� B��
��|���fa��#M�y@0�	�K�Y���w A B?�T���v�F<�K�$6��=�@:@�	V��o%D�o|r�ѡC�e��vww1�E�iǓVj;<=���w<�` lQA4�i�� iR���2�kά�N�"ů	�ϧy�Q�')�]{��'r��{��/�o����8e}����,C��ׯ�}�x�ė^'�k ��O"s��Q!����?��p0�z�G̬�F�b�!��捛���(�}�Rĺ��E����>?��cb�xHP���4d1Z#Djӛ1�� ��� 
*d��i��h���ܖ��/Y��� Jd�Z�^�J_gy1�O�OC���75̌$�VO��tc]t{����1
�B �� �Nr������DS��|�9���ٰ*����/�����_��{�����R���ܛe������Je����anXB��V�L�.ݤ�}�k���/'�����"��&��K7�����^f���l�|RM/���>���d��;��t�kr"b�I����Ͻ��7����6��c�i��^��ۛ�9礎H �Ci��	���pN��+A�����o�e#+�z=(V �'�@!���H�5 Cf��
�DP�i����K�C�Z��i�_`��}�O;V�^�Β ^��|�p.@��Ĕ�<u���ܔXͲ^Rh���a�;�]"�)�*�7��?�I����[��9��~�s_:7����)�YGH`�� *]�w�p���?V�S����W���N)H�3I�TJ�g����>�v���x"��>u��g�(�>92Y��U���gG�Q�^.���P'����R�͓��0V�Ƙcjͽ�[�J��������8�<D<z�>|){�� �d�<�)q:<\<�`f���wr�@��QH��
|q�;�?��F>2sC�S�ӌ�A)���p/�[� J��×��>e��$��
1T���DT26:)4kd���V�@`o�W��2ɏ��k�Ի�V��W��g��P�������vP��4���f����C2 r/;?�hP��I����1Ed�[����={��IZxo�d2��Yi�t�w����;���GH����؟������"�{�h��*Vױ_�'+�W�ui-m-��b�r�#�p��<����&�1a��~~CSt�/���ʗ:%!"����D�Jڃ��o9sx7t�p4�s�C�Z��&�{�9�4i���q�� A< q�}�$ H�$9�Oi)5#�T��Q!��M+WlV���{�>��}��
�4*Y������ �2L}�x�2T*ػi�6�֥�W�+�[���p)B~2�j�?Q&aEdX�`�ɴ?����&��I����s��ō7�Ĵ+���y��\�?��m��3� �<����X����8{�,�y�\�y�|�<�r���w�܄1�Q�݈/����')�ە��+�< �k#8 ����Ȥ����СP�#�w/F �F�>��H_�^��\ 3��Q�0 �p��H�N���'ȳM�g:'��wΏ��=���Ɣ}3�� <�T�J��t���e@B�����Q�"�(HP�(S��?��2ڔ�ZUي�D�����Z0�MgG����V5+N��~��5vww!lmmaV��Y�&g�v.<���ڤ�6�z�hU� ������/��,��;��;�i�,�2%�u Gb�s6�<���!tu�g B�����D)�{�����Y���f�CT��t6���;�B �}�[�����5	}(���q��*O�.�N������Qณ���;<
����ó޷��]�J?h"{�`�Ƈo���so6����G���g�I��$q�ϒ�F'�}�[>���r���R��|�����}��خ3��ѼDf>-)?7�z����;�=��,Ͳ�F�C��J�� �B$"�
y�� � �uI����"D*(f��U@(��(&<	^i�"$��6+�B͊Ib�*#���H�Ib�!,���Դ* �\� �Z���Q��ڷ~���ج�1KD�̤�Zk=�I��,˰s�^���{�Lo�D����?�'��]���硲E���Rʧ�F��P���]���1�J A)�s�Cu�N��h��H�E�[աýx��?�XMY�:�P�^)�%L��"�A$�.H���A	)�B�7Q^�"@��h&�'��{OeY(�*��!��@/IRff�C<�V�v}�=��s�����G�^������ɓ��f���G:W��s�s�F��Ȳ30Z�9綈����.z����k��@�b��HN"���&�1������2���N��C���T�:tx���W׈}\+�t8�`"�s�9�e-.X[�;cHi�+�b�����;� >8�(xq"�A�V!��"B�YvΒ��O�S
���>h@3k��QJi���r�:�U4~xk�׽D���y>��%���eΜ�A�g�u�&�b�Clll�V��t�;w� �{���]�L�iVLo�?�?�ү�گ�����Y�)}�lr�f��mKfa�%�HH@�P���k���Z�[A��o]"���P/2z`�(m���Q�yo?f^R�����q�w���=���e�b D��B U��Xc�R��*Q"bD�/>HHB� A�D%�+k��W� +"�	�FR313)�t��e]�˺���b���K�}f/�Om����~���-dY���0�L����Z��
E�������o~3�~���Ʃ�-�������U���c]ҮÓ����Z��A�RXA'�����f���6�� "D�s�p|�:��p����C��6ډ��$ċ��z�ZnȐH�'B���\� 9 �&�q�ИN���i��b0��H O�!fM�}`kmduPꕣ-/ū
ߊbȂe�W�o��hI�ॗ����3��bVL���I�N��:�1
��֖ ��Q�=E�� p����_�tx���>}�;���Z� �L��D���L"� @���]T�����^Glj���*�{����ѣ�� �(����v���x����:Q��*}ǭۼ�>��<*�)��ޤM��"���dfx?.�:�13����i�I��:Q�;����V�ݼq�{�(�,� C�9sÍ>f��s��eQ!� �ij��A$yֻ�on������S������H�]f�ƀ��BbK ����zi���0F�V�4�6s,G_�:���Щ}:,���I�����!e-���z�!���2�h]Oo��kq.j�I[J�<�\�&� �M�D������S��E�/�p���}!,����^�G?�Q�>s����-����j_��V�$�h�&߶3��s�_��_�8^0<�;U���p`�@���wU�6D+�*Q��(Fb�# �߹���Б��G7�u�P����Y�t���f�ZYRט�ԫӴ�a����ץ4Rjq����Mۦe"��UU+h�s��]�~8�{0�ϑ�9^{�5|򓟄��,K�z=dY�;��6��eY �4y���*���a���W���~�N��/�������rG@v3���l2�['N�����c�q�rVS=�L�&AE��)�$���CQ�0f���:���YO���,���]m���y���GᨴG��[���A���<i�`y]*�G���qT��z><H�����쿣�J"�8�����p���W�պH�"V��8LZ�|�^�m>h�i�u��u�~�w��yy)�М|�Fa���������.�3`{{���'�$��[��N�:�O�=�d��O�������+ ��#|/��F��W_��ߟwtFw��ǟ��'gI����I�M�1���ꢬ��@�A���P�S�^�`�F��u�p0����A[�jGyv}�p� m�|9���"ǘ��1�ͺ1�<I�4�x<FQx問೟�,^}�"���
�~����p��M|���&�n���pk�Iʋ��w���_}�T��S�zU��׿n�^��Q��J���Y�5��ΖU1T�9I�*ɒ���&676�@��$�,�+��l���Y���?�>��C�Ԣ�9�A��p(��~{��6-��kCD�A��Df I4�"xo��p��ŋ���ckk!�z�y�<�#�{`����0�_*Q����n}�W�W���_������Lっw`���K(|;�^e�NΊY��e���I��Ι�8��^�\�qeY@)�T^p�r ]����z=��t<�ѣG�i��������|���w��1��qǿ�$�q�A���D��t�T��/MS�Ԧ����㻿����k���ad�<yŬBUY��E�߇��wG�����ɫ�;= �_����#�P�g�;5���'/��3+���~K��D�S���p!����>qr���Š߳��P��$�;�M'��"(X��=�*=ݓ�QX���t��}ʎ����3�(p�>k�O���,���I��У/�1�����>}�}������_��!��41M.�9�#��R��z��{8{�,>�����q���:����O�<	[9��3L�%��iT��wn��	�N��?���<Ҋtx���J� �dU��
W��/�$����_*f��^B�C�~n@Ӽ׳y��T�M^���B��#�S��v���Ӎ���G{�����yW��t�5�>(b�~���j���+}O����s�~��7/��(�,K�$	N�>�4Mq��&Ο?��/�ĉ �z=�GwB����: @�|�]��Z�����v��V��3�V� ���a*
C��>#���~os��^���Ui�W�$K|pN)�$���{���F��,ଅ��������ĕ��Mz�U��;��xԤ�Q�q��G���Z�8��o>z��1���?�wl?��w����~�m�z�u��A<Z366�8u�Μ9����x饳x饗����(ב��Z��ޞ�����1�ͤ��{U1����tK�u�궹z����f�u���KL��`�����])ڝ3"٪`�[;'w_��˷.����ڀQ�0����1��?�N���#��;��?G��q�5MSlnn⥗^��/�������`���[����{�5��)��@��ۓ$�RUe��J��i�X+����
� ��}�k��o���1�L&��A~{�u�����~p���������);33܉���IY$voJi�(�f���z!�JA��^����&��8�E&�A��񷸬�q�\wIBz�N���#\!����*���8��0��m�0_zx���܌"���:y�Į����L��`�.b2.���9ݻ��r���Ǆ�1--}��k�5eZ�?� (Z^��}|��,�g��Z���o;��#/�9�bu�����f[X^�`������i�X�+����o�w��ς����P�˺O�:�q��n���s����X)8���[*C<G\ybu\4�,�=��j~�����b�7k˥v_���a9G\���2O���i�a���v���	/ƈѦ3Dc�=�b�Z/�)��$3�97Oc�X2��p9��u�=�ݞ�_�� $	��:�X���`���^�Ͷ�9L�S����g�;}����!@��߁swo����;w��w���K�� r�����ކ���wn!�����7��ڿ����� }s�G>r#��>&����'v:�}��Ib�щ�TU���$Ku���ΓىS'�k�����[��;{�����H�(�.ԄB��-� GY�c�+ R$�x�ѫ�iy��ݣH�Q�����p��I;~_L��'�-�b����v��U�О��ui�#N8���`��UR����#��d0֩MW��&KXS����H-ױٳ��X�4����q�:Z�i�����'B�4�,��]�vߵ��>^麜���O�6��y������m]>��A$pRH͵��PUJ��9"Yr��2���r�:�T"�l6��I�W�r P���>\��Ƙf��v����kκ����H��X�Д�Y7c6���hD���oږ��c������6Z��<�Q�2'ζ�^݆59�~1fBX?�e�܂<���ً�ؼ|����곤��]��n�Y1��.q �e	�666���1�q��-h�������&v�<��    IDATv^�Ω���
�{cTU��~�����>�*XW"MS���e	�1�2���&|��݅s3����W�^�z�õ����a���i��+Z�[Je}R��U�4K�,K1&U�1��z`����o��y��M�g�z.���u�>�Y�b ���y �����	��t{�<G�"<���(�������Ԋr�S�:��������-�����:�����_|�o?�Wϵ��V")\/�	��}���M�"'���'����j�����
q�5�)�q���o�]�u���uM�޳�j�����:�6n+AD�(2qR�u���*Xk�$YCļ�ͲWq�6���eu�c��Q-�uH��9o[-��QJ�Z�(j�,�:���&6u,��F!���4M�k�[%=�ǵ���^��4MQ�%��+�r�R����W�U%�M���^%�]���.�s���?��mߧ�~���ƶ�Jg��C�����F���}�6nܸ�,�p��Yl�z�?^����Ac6��UƧ>�=x���B��_�1��0Q]g��G�L�(�+���c_�/_�r��O��>�?�]G�{��o��ܻ~H�4���$�����_����Y�J�P�4�3d���i�ʻ���$�~�����y�����G`�B A 0Dh!'��Ȃ�3/���C+u��v�x$ȡv��S�����C�C��=����X�.�0����ww�q�W a��|��U�\:��~���)_�:��z��X:_�	#�����C�˽�������^���������th��D��G�������3N��2ah����{�Z��������2��%"`�8vՌ�&>��B�{����@UUK�_]�UHD��)�2��<�6̲���&�J)h��Hk�L�~Q��n�+n/�r-Q��&�^:.֯m���5�Z����`�d
o�z�s���kױ����n�����S헠uc���^�V�G�g��g,@�[��v�m���R��~s�i�$�%�~��e���1�
a6��Zcju��*��H����}{��)�Α�H��Z����PFa4�C�ll `m���eU�t~oT��N�������]�rep�ʕ������w#�c��YQ|S��|Wk��^oP�keU��ͼcDBe+�����i��=,��2��
��1X1���� ��C�jӮ GġESp�[�:v��y|8�'���k>��$�i�A�r�vB��a�')�`���^<H����O�,�@,@ K@@ I�]���(���� �

Pj�vi�������b�W2(���Z,߽���O��������ʣ����Y#MR6p������= ͏����ܨ�/J���6ɉ ���.�H� W�Wz�\��=��:�*m���*��H��9vU��][�i��/~��#�J^Y��$�L��,��i���ܼ-V3/O�(��h�����KkmC�$iHO���~�~��,K8�`�bY�$I�r��G��LTۤ�.B�e�<�ֺ���~�'��J� Sm�����jz���{��������n�����)m�3�IDP�e���y�<�e��Z�5i�ĭ�OJ)�8qb��3^#�����%��_$���J)8琦9�,C0��*��N���� h4 �n�� ;;;�o��B��{{�U��V(K����7�����?�?_��?��3W~�J��u8K� \�tI�<��Zo���`#1C����D��%ȧ��,K%5�1������&�u{�w�ڻ��n��hei�� ��H�A��U�C˳������ e=6i��P���ں}�(���G�i��ïϭ��dd�\m��uXU����u��u��:����Y�t�գ���quP9��V��^�7��J�	��*Eј�V���sr��t��a�'�֪p��N	)��2�V���:ڪu��M��HE��d��H�VդU��n�6I0Ơ,KE��O,�lV�إi�,��~o��\�d��Z'�WPS{�KhaN���sB �f�z�}h��,g(�
֖71� B�N��sq~=�*$I�$� �9�RcR������) !Ծ�����'���5��ޣ,K��(����Hh�ב������8����'c�y���m����j�|-�tF"I�Rf���9�b&�K�d�'ܐ�<���a��Y[5��K�m�m���	���}3�"�t�5�3�e��aC򫪪I>���y���w���7Bo���g���y�&n߽��(`�T�w����A�o�������_)�\��[W��ӻ�@:��PIP���3��l03'M��։V��}�W���<K��r.��i/�43 e��8�v�;��w����=�2�I� F�F3/���Q�*�Q��ㄠ��2�}|������"�>�?�|G��z�<h.7�N�h>�������7��'���Ѫ?�:��J�ڦ��b�6�����b����?P����0����^����>�ܹ��h��H�&4͹ԲIk����fR^%�"�4S�
���U��6�j�'N��l����T��6o�rEu�MҢ�U�H6"��L&�m������ �nUU�iq0`8΃K����F4�NU�V�r(60�Bb2$��V��BeKx`]	g������E9�b�43�����3i8W�*\�`t
m����MK�`a�<u+�I�Um�$�_
˪� ��su ��<�/<�C��G�1޳Z�#P% ��h9� ��i���~T(��h������Z�,� |�͘Q+A@��*��j�Z���.�����X��A�1��<�c�Q?�����ss�n嶙����gM����m3'�u��֪��c��������t�ɴ�d2���&�Ҽ���mܹ�k+y�����`��~�O�/~��~nt�C�C���I_<�������O���W�~f�+x��!ȧ}e_~��A9����:�]A������}�=��aooB\��5~}��F���aJ�B��Z��P��}�v�O\�T�'O'=G�(��0�t?8�x}��YM����S�$�e��k�LŴ��iژ�bPF|��f���Gr����|I9l�mSO�H�	b��_"k��ŋ"��<jD����qRUJ��YS�U2֮�AJ�`�[�O������گM�������?˲l�Ik<gUU͟���`���~��O�UUa:�b:�6�9�&)'N�X2oF�e5�&��H6b����`{L���n�]����Idiִ�BiT�/>��Q��D��c6�-)�JŔ/u4�IL��&��s�9�9)��Y)ds����x	2'm����$s���n�f������Q�Fǀ�,��=�R & ���ʞֵK���KY���sEQ��k�8c@2�Q��8�G�@X(�޻:�̼O���b�<��4m^ʪ�p0��j��E��e�,�1>/b�͊1��:TU�J+mS���צ^ ��_Y���Y�������Y����ǰ��N�;ބ�B�����2��5��+��g����>D;tX��"} �˗/��D��>m�R�n��}��R�7�?jg�~���y���i��F�Ėnp����ƍ박ŭ�w0�`t
cR� �a��h�m��ќQ��'0F`��U��c<n�S)��1�ALC�����SќI�RY��H�=�B���n5o��r����f�iO�q"��/�!��=�k��o|�����b�g�T4�O��`6�5���(�E$8q�h�h�����v�^u$oO���%B�$	��>Ҵ�o�6FD�B���&�<�s�Q�vvv@D�lM,�/Sl��O$h��i�6�p8���.��h&���Փ4M�RUU=���7f��p�`L=���]���X�����4M�mj���� x���`&��cL������ʲ|~�rZ�����B��&�跴��ь���Y��r�ǣ���|E����Z~\2W^� �^��c���e�2�n�:[�c�/����{Hu=>!��=�E�F�Ў�m�x�R�y��o1��DP���CL�R���ǘH�3�&��eH�UY�:���<R�ZL�$&i귪�:��$�ι)�&����xi���\��u�������9�<���	��s�u>�P�~�ߐ0V�o���
A��?h},"��A "�����O�⠈-)� �>Q�E�v�(TUiʪ�B���AC�� @���QPJ��B�i�".�(��t[�V� ��%`�"h4�U &��V�����?��~.�O�. ���Ν�鷾�.��r��+��x:�_ �M<��}g����/�ߡ�x��/^��_�rz��;����`��OhCQn�E":����r���Z��t�1͒�x�U�0OQ��Y��x��N0�0)h�@`�5�Q���	 +��	L�!XW�*-�^V+���<$� ��P���i�7�j�@[-h+�A���1�����;$f��,�1?�z�F��>Ey�7�0^?��C�e9Z5q�	fkk�1_E�,��#�&����s��lS�?����S$s1:��NTVΕ�5�iH�s��%I�y^����	3*M1��s��h������M��bT��|T��m'�8�Gu=/�}!���X��9�D��M-�M������*g����TB���OE��&+����T�t�U4�IӶ렍��,ʲ�u��'��/�[�H{ۗ/��2˶�p��+�;�2�Ib�D�67�y�a�J^$V����aE��"��W.��]z���lU�HA)��F����0�`���#��|=�����C�j�"�B�9�����_<��������ypZ��jk����ֆAP�}]��Kkh�ʲ�1	B��y"q�	�X�֋��Ԗ'�� !	B�P���&ˊ"DD���@$�a9�IZ�Ê�3��z@>t�\����xϹ��x 4��$}+R�BX�E�,�$RJQ����2O K �CL��9��'�@`""�P�EH <�aR ���zAsP�,+vD��k�l! $̐���$��I��;@"A��B">!b�U�+b��Y��_��	#d��UT��t����ݟ��y>���?�L����A�  �/_N�a��]�PN��O���*����dF��aY���a�;߳�K�,�$�Nz�0��BH����N�X�QUD�(�i�<O6cR� B����ij�ۊ^�,��A�h�icTs�Z1\�����تI�p8�p8D�e9��"����⧔�x<�p8D����d2i�^���<:����l6����� ��d>��n^��R��ͣ����s��\�:|��R����a�##�"M3��1�ჯ#���H �4C�&K�l0)H��6�B�#&dUK�.��AԘ�j�!����è�(�k3�yZ�������o㱝#��j[��8��<k �s��E�uDg�Ӹ � ��R�pE�)��lND#q��D9��s�U��¼��m�w�?S��ڼ��^ӿ�����IUU��!oT�73; ,�T)^'�+�l�JIT�j�#�I���/�H2�@��+"��M~��פO� "�+�zH�E��9�HC)��0����yP�dA�h�l]pD��5�@��H�/����L�&B^���y�l!^+dV����}W@,
�"u�w�y�uU��^o���nN�4���LJD�H@�S� �'"$@��Je-��*[��2-�����	@��J��r�tU@��HB�E�D��G�1���H $�A�AAI @������2 ���sW,AẀx�V|W@=fQB<��D��$x�����)	 1	D��f"�~�pD` 3�ibė�kbH^)eCDLM�������(2b�)E�$�'&H1Dd"H�2�� U�{K�f���Ay	��#;�wn��N7�����L���G60��ߴ �ʕ+-/�>��7��{��{�0εҼٓ�U����T��,M�D�t��̺��?���;�ub��^� M�4�$�xv�Bو�H��677[*��RSTc�!�m,"jT�����Of�[2��sE�0�����H��&f����*���P�A��2J��%�|���H���KD�Ρ�*�������D�Jկ�<w쟓�:��CzC�S:4�~B��O$ޕH��A��{("�୅���5Rc�ZCs��! I3���ے$�u����{ddfݺ�MQFR�L����ؼ���K��z�٘���Jf$!U7Ш��k�����<����F�6���~9~��s����:�k,�U��)i	��{kG�UCeA0���9X� T�bɵ��&$3�8>�Ja%�2b�,_��^ � n�w�5в���-^�V�(�c�r �����Xs��3� ���{@+e:^gS��cV	���%�@�(ux�Zz���������ܘ���P[�}fh$����C��df$�0zD$]\\�܋��{I� `�,�ٶȔ��ڳz��<"Aw7���� ia�7my`�̨��XI���ԡ��Q3��Zދp�ʵ�#	�^m�������$ #@3/f�$�H��+uiXҸJb*I���c����X� 
@���5��v���2�e$�$4��w ʁ]2�sl�"C�Z)H������&�d$W	��=�Rmm	�F�E���g��$�@l�F	� pA}>��/ R�(���W�JZ�4��\�'$I�z-�nM�[�f)K'�p'�F2�S* D1 ����ک�m%xEr���&��##/(�'��mD��v&܂hi6��2q��%6 ��-�-V��kt2E��EDTAFh��b�w�j����=i+i"�vfv'��H�+�Y�h�����>��s���m������=�����������������O����T�e�9x�ʟn�G�/ß�c�'�0���l{r���N��R�����0_G}�a���uj鬐����k$2���� ��������G'���������]��a��~z��&6<H����<ߧ�: 뚫u] �#=߽��>������S�=J�?�ൃ�^ŷ�4Tv���NN6�˕�7N2�`�۲f�^(�nΖ�S	'n��ܐh	��B
�XriZ�h�i�D�� ��2-
����ѐD�	�U)�Ī�(Kw�4YA��&W��2B-!+0�2E��.3�����s F�$��2	�18��~��Ps:�fT�L��*�#�be)d��0���`BA�a����v���PI�̤����T�

4)�L��f㍹M]H�$P�)d��L/t/���%Pf�D���%�$#��,�~��\�2QA�R�^��(QS�H+���֖u2c�֧��@�P���}D��RH �G�	�_� 
JI��!#���:=Y n���}�v���Ğ�
��d鳼1"rE`�TI�)�h-/I��l�@b�
Ҁ0�М3cf���A ��2@ �4���3��h��o3�k*�F�SP����#���f��I�+tC/���u����+�@fJ���L)�H���QIb�q$A;%WAň!%8�;A'�m��  ��J��_)�KȾU�^���NED�7	�X�k +�'�8�l����=I'���6�k
��4'�Hy �m"�A��ɜ� ��p-��M�yVk��T#���nU �������ni �B��|&F�% M�`Or��IR��%��?북_��~�ܜ��'O������8��c�>���իW�����G���N�yi�+���"�|���T��t7e�Z�l�O`�֩�@�2ġ����x9�O���qdɎ�s>AB�p�Bz�f"p�jzT��ʠݛ�>�a���M��B�h�;�6��8s�������t�?4�P�5��.�D���H+�Yk)���$��Q��3�\���H){>O�{�ہ�."=�v �Q��)$�v�9�6�	 ��F�aZ铨g��Y�3����0M�v�XB2t�8����L;��׵���Ief�gt�X)����������}vP3�sg�jdP�Q�%47[����1�B]�Y{>-S�'�  �IDATϻ� �2R�y��Պ���80:<|�gEĆ]`�#���fB�}R �IY�$.��P ��́��X[�� 2W�Q	,��8Q$Ԛ��_�֚�e���fՌ�nT��[�sR�ݥԤ8egD 1��"A�1��,)A������3,(JU�$o�>$��=2�Hj{�5�M����Ho� �a��!�*�$�9�	��-�;�/��OI�SZ	��䒉;%�ILNlEn��H�S3���]n3󝄕�		�TK�#һ)H6�n���Dx���^]j��!͈�Ɔ�J�(ak�H����"?��-3�B�h Q%��ߴ��ɖ�7� �L���r�\�]�E�B�Uٞtɥ"3P%x,�=��@��V⍓�('U��q�d�RH����+��{����Lc"E��\͆�\���U�G08����6Rq5�F�3$�L�-�&���*�+w4)���IM��t�w�ߺ#����$2�-���5�朴pG��(�� k-�k�gt�TgH3����Ӭq���f���&NOO�f�������_��o��W�^�v;��x���g}@�Ꝧi�L_���6?����/�C/+��n����M@������8��$Ǻ)uܞ�T��m;h,�����=�8�����ﰎ���x��#�Ɍ#���*/�;�΁G �R��(�`5ph;#C���PD�A-"��A�:�$W7��-��Ks�=���*)�fls�w��T�c囓M`-^n���m$�������m�k��[@��F"�|]��B2(�P�d��3�b�������ڕEY�|�wo�͙���s��O?W�g@:�4Zs�5�W������L܁E�H- �N��WI)E�Ҋ�eY���.J�p۠���!` 8+u����	��n [6�͔�kk�����( ���x5)��x#q6b�Y"e,�˺�wo���,<!yzD����~�����ȑ�9����ImP�+	; ��!'�čB3L����aߦ�Nfb/a!1H�i�:�`�"�k�)�f0/��~��Z���'f��r�S�l0�Q��s O��g����T~f�gF�0�.�k�R�\��݀�!ٔZ�^Hy��i����e���� .����f5	�������ߍ�˔�ؙ1$EH�D
L-���vR����H��B�!�s	{$/�!I5�A�.�?P h�0K��( '$nIJ�(J$�0H��n�_"4���쓐S�D�<S�U�Ud �A@��um��+���\H*"7f~����R*;;�R�LH�6������d�_|�/hȬh�$Z��R0�h ,��KDld\���v�kF��b�j�Q�eb|)Е���
V4d{Lyr�zY���� r���8��` �%w�1ǛKRb���ZaZ��5
IX+���4�P_Yï2��L{W+�Rָ����zJ��lssz���;ȯ��*�����=�w�ޭ_}����k�믾�˯��C_8]�����_���o�����������_�ի�����-��|����EU��,��Z��0�i�4����8�G�mj����A�r"Pͬ���D�ѕ �g���, ~H�t	��;i($�~�F��9�\�eCGx7� �M�i.���  G%52Iq��ݲ\oo�-3��:b�1��p�S�F#�&��*����\�y/7F�N����IO133it4�\D���)!�{�M 2%3���fZ�"��г��֊�p�EȚ絖��g���\� ;�� ��s#��0���?���[Y��; 3L���\��d��-:��.h�0)���7����D~"� `�]�R#�~a��M�|
�3 ��ncm����	����w�~���1��k�3|������ߓ� ��ไ3
��wmk��.)�q߱%�g����i��c^�<!��]&tA����[C���F��F�fƧ��<Д���_�"��(��� |�@�X  �[%6N�*�6�.�$h� �=]��,�3 �J���[#/	m�)��4�)��ĵ�Sx�^{P%�;�{�F	���m�.�ې(i�-0p� �� }���L��4dg^nL����܆�"�&����r͑կ�r�(&��y��%�;I7�o�	if����\R��D3�-+�%z� '@[4��#y��}E�ȬP���wsY��G�Ӣz��f.w�����Z Jq钭A`�{� @�=؈@9� 9e� d:k�{[@k!��� �sRՒ3
��C��Y���-�e:��<���V�/(xZ��F,c�=��Xչ�7f*)T�eڍ��L|6���ʥ*��lD�(k��������>�Э����͛�>xSk\����Zk��� �Ln�Z��,w���`!� �Oc�ئi����NNv����z��J��>׻��ś/�͗��իW�c�������} �ӟ�����nj�'������l*�_M�|�����?+�gn^H�����͆�1���Jq7�.����5���I��3�� ��@�vR��� *�VX%5��A��4)�̱��W;�+׌Ʉz֘G/+	2�F�5���ܴ�g��ˌ8����R:3c�|ۢ���)�Y�&h t�n�ì������V�$9�B��.�fU�W7��Z��P�@��:��eYwkks��9i3�k���^~'e4(�	��כ�Dg$�م�B�R�m��	If�
�Kwvyf�8%���N`lۥtr�� �EK�]223�Pb��zrL2���R˥�C�ŀ�T.���v��D~"�ԀJC�~)7�)u�J��h��%]��IFP��Ab�sr�����$]>��� 3䚀���� ��Ժ��^�|U�%8#1��B��̼7)�N���a�zuHK�c�dy�	��.�*��	W����Z �t�@k0yxfJit }�?�?l��g 0v�%ݍRKX~fBK��akB�H	)�M��Q�Z��_����B܃��F�P&ҽ�݅�ѫ�#Jos���M��R6���um�R�ko+9M�L�<��@����k}��w�����e�p��_ʬRF��MS���� ��d���q�I�vw�ֺnطO��|�u��~��N����z2 �ݨ�:�o?��D%BelH�-����C������,�M �>��0WL��^�]U���YK���sؕ��~�eZƉ�ɾ�����%�' �a��4ޞ�v����[�8��
 �6��n�?�=����˟<�����ܞ�ɓg�!߼�B_~��^��J/_~�������c<�s�AAЭ\���FI�M��fu�/	~2��8����?+4V>#����W��҉f�&���TƗƣP;$n(�ӱ5b��LI����7�HQ`V/�(R *�eu��g����dH�h&5>K��id��t�����
3��NK	��B�����
p��0W�S�߈�4�M�U H����m�� \�-�u���J����q;όZ��kD\R�IF�>y��-���Z!5��D*$:��)0� @E�3�mf�+RA���$M�}s[{i%uH�5E&��x� 3����DO�Q�" `�`�,�0�JQf�J���
q%R;�H{ �������$��0��0i&	���̔��y�����L�d�(�/#��.����.-���(�@���i��?����Z���³�x�̜N׃֨�r`g#��l�ZoKQ!}<XY`YZ��eo-�����E���a ��{���,�e9M0��Y}y�o;��'����uX+[��� \�8p]g�:>Lo0σ��;��p]��6��eYUʠy^u�G뺰��q\8ϫ��է�O�5 ,֥!.�fX�}[�ۍ?8��k?����у��:}��|�߾̇��>^qh��ǫu�a�t{ sð�_�,���3w�u/,}�����q\�����_���z��<m�������.���۫~-oa�ߟf٬3�s��f�A�����(Ĳm������ v��w��x��W?xN/_~}��ի���6� �1��?8��W�����o���nv�� `:�k��,���3񒴉�k�Of�A�_�`@R֋1��=L/�Lu��ƍQ/H���{�P�&�)�\�͸d�dC��� �������U�p?�Y$VB�LUR��AO?1�i�ש|����h��{ !r0 �v�c���4ebDv�����(����1���=]�v��,LLh�AQ$Y�7�|XVZ63Xʰ����_m�h����|5++�A�d>e�T�<3��ߊ+���d+��%�V@rgƝ�-i��ꆖ�Fz�֙(��,ꂺ"�6�`fm�0��j�)V_�դ��=f#
V���'w�hfvkV@������fV#su	�Ze�ȭ�uW�����꺟5�Z�=�N#����6�~Ts�Ojp�c2�NO�ED��:�v�SEo�>׋����o���>\w\���;}��x��+�˗_�͛/���� 8nw\����a�����_����V p~��wi���i����xr�A�<�	<�8���7�{NS_/1�a���S��ސ��Jv��ZƱ��c�����wG 8Y>�P�f�q7�=:�o�z`7��$�ۉ�2r��sYfN��;��$���fk��i��z���V纹)yz����������|�m?γgo���}�;��O?}��	h~�K���ׁ��?�^�ze���ן�>��9�����5��_�����_���Y���>���1�)����c��V��4�7c7>}��_��!�3酴�3.���XO�� %�ޘC0 TB'�vNh��7���[*�tG�^����L��>�N�>�&F��pD&�P���mY��g���,׶<s��B�+ɯK��� ��xY����\�J#'4ݑXH�\[�@�j�[3�0r=T�Z�Յ�ȴ-����P�����9�8	��3|=d��^�e���ζ�"���
��b��a��E���R�KQ)m�`�9Pb]�܋�|�2oUc�[����<�P�ڙ��� �8�pW
��K,�iXі�2�h��ke����9�$����\d5n�Ǫ�o�Lӓ��g�a��cĊ���E;?ǰߣ��5����\Ob�R�6Sm�5y9_\<���Rʙٮ����N?\��!�t O_�9�ޯ?=,��^
���k�3#o�>���#�:h�7o�����_~������a[�3'�u��x/_~͇�>\��s=�{m��7��9�`��/�!^~�/.��˗_��GV���ա/� �1��4����O^ճ�����~:n��$_��!����2]��O;��Mf�@�!qE`1+����^�]| �J����N�v�׊�V�j�½�k�rH��)��c.<JA�>V3���<�}�2r&=��x+"[]��W��*��e.�e�(�ԝ�<_m�mm�4�-��,eЪv>Ȃ6S��tW�ڗEcC)�J'�9xk�9֕��4u��a�0�˲�f�����Z���C��I�]����q�����,�L;%�%�\{?����9PV2^�Xݹ������n��2&�I �d���6��%6��X�^e�s4�~�+e_���f����,���F������v�Dggo��_�;�����<����}��>\��I���#�x��x��x��o���> ҽ[��ۡ0W/n���h+[8�+q��iC��Zc�CT.�ʗ���G�0���B����S>%=2s��P�P<5(s�b��t�iLN�g��+�Ĝ�����Z�s[�7m��c�
 eַ1�S�=���|�7�� ���0����nW[[��C�J���t_jD��Ϙ�%:��o ���M��#�u7jwW�r��"�g�%�m��ۃ��+Ǯ!��>��`��lnm���!��A� gg�����_�`��__�_�I����<���x��x����s�Q��C�?�i��ؖir��l��"���Ɓe�lM��>�q��u�6 �����ף 9[���ib���RV�y��\� ��]�W��Y�Png-ۑ�Ǝ1�4H��q�C��~ G��t���@tqq����_<�A�c ��{�ꌞ=����~��y�+ �?}���<Ԁ�P|���ݴ>���1�1�1�̠�a�'?��}��%?}�������/~L|~�����ы.>{�#ktd��/���x�� �~&����~3XzD�����������B��K��    IEND�B`�PK   �R�T��!�D�  Ԟ  /   images/cf2dd1a8-295d-437f-92b8-7fcc138ae9be.png4�uTT]Ň��z�iF���n���n���)���fH���|k�e��̜{������މRQ��zM�a��J�?c��4�<u��Ar�b^�+]޹��<�B{�������\�K�B�EБZQq��SH�y����87�����o����b_�,��9X]�'�O!_�YM�cMO�S�ր���nS�[#~'���SB{��7���	"ݚ�g��)L ŪU4y�����[h! d޽�v�YHl��T|�S�F�>,��	�Qr�4Y�@>�T`Kc򆓓3�����=<�$$$�?�dff�°Ȧm�A�\W4�^l��r��!S%u��m�=�-Uv�q���)$%�_k8���恢�u�����G�j!��A�(g��r/���n���OOO��\�H�ژW��}���!�A���b�ԟ�! �0�,~*<V�i$o���=_���YD!�rL�ӶyV6�y�Q��>�K;�MV�+v�3�0-���c'1�] %x��8��������.F�6N�6�j����N����L��z���D�u�����ဂ�Kh�#�R������۴Ϝ����Q�J�w5�'�TB�G�琄����q��|����ٞ\9�s�\Ԟ���A�AEA��s ��Z5���͟���<s�P��I�̋�ƥT3�Xq���fFZ��d�F�h錓��Y]����A��ur�bR�n�쐝(�0X<(a#���Ό��Zg30�2dq���ai֭��N�\B�p��n���M�ɴj��$"Tޥs@�a}���(�B�3�����@T䘘����gs�@?J+�&�4��@~a.��au��E6���"�s���s���-���u�n���b�g3d����L@z���L�͑�숀r�{��͇5ua��p�����52�)���~I�ό��N�x~,����TI$qɁm���>��,�4��_:��8Ej,�nT,�"�dr�3���zmj��(>�>5Z�7�}KK��,��y��U}�8�d�ݝC	?�3U�9�O��}&��̬,1�n4J�Ŧ 
`	uk���%��#Ȟg�� q3�(Q��> -q�:���Gq���9����A`��QG,.I&���Y��I@b�����]鶟W~^
��a�����O�	�镏�~��2Ţ��;��������/}���;\���-8f��v���0���������U�4�;d�U���h�OK����L�/݈_��)N�"�'��!N��sFr���i)�i9���I@�@���5�8�ۈ�|*;	ѝ`0M*hڂ�PNX������M�Is���N�����a}�������ڞ�(�����`�5���X��هl|��2v���N�feC
R靾,�X�d���b�J�>A``�����Q�F��=)f5�������kd�3?*|c�3��!��(d�(d���Y�"c��2�����W3N�+�Ӻ��􆇯�)WZ2��حwSt�n�`��
��u�&)W�a5/�#�� �xз���۴ח�_!��y�g)�n�������GC�I��qԨy?�ZS�WB�R�ꝓ$�{!X�.��:F�!nn��Pξ�Gbl$V��+����N}��N}_�P_��Ȩ66{�ZO6�W���J�GMmm_�I#��ˤ,UJ�W/b�I�YRx��~UG�u_�6���,�wan�ɔ�2jŢC��D(O���;]$!���Or3��.u9�./���=�[��u�^'-�6T��D�?�x~��H�/;;j���5�R,M��ݵ/�	2����"7�掆�G�M��}gI�j���1m�l������m�#����|��K S��JJ����tV�fqZ��f��<{�x�{�o�D.%k��76�Ag�LD1_Y0�ˋ�j�eP�8GCVqY�0�!�o��o��9��d(����YU�s]�tY�~üxB+o��U'~(<}8��zN�\�a���1
�ơ\l�_���4��N0�Z��p_-Y��Oe�m�/}��2L��6e�N������}7�|�v1�m&խC��|0��EI>�"�j�6u3�B�[��p��� ��F�G��AB��w80@�^K��;�Z�g�K��_n�$ɾ�qӭ��1i���������$HL։�� �#�,2F�F�	$�8CB@���ʧ*�q���G{j2L�UZ'A�����ۏ��=��m���Ï
�o�>�XB�����q��k��K�h��e�`�aэ�ܲ�3�` =�� �"��օ��������T�lwq��T�l�,.��h��樻,�?>�?Q1���Ԙ J�bvjD���i	�$�������Ӓy[�4y9��Ye�����
����nad���;o�(80qF��� :�c�ǁ�YN"7�ƣ���o*�ߚ��"EyQ07�=�Gb͏�dc�g�3��gB'�LJ�K������W���͚�46
&��H�Dwp�}���R��{+<����,9������݆W?>��p	�š\4BH�C�83�#�\�a(fP�8t')O�3Fn�t�����n�H;.|�uE�P*ư�v�Wn#CV}�PoΩ�	Ҫ7dm ?��"��4����yV��ʊ�$UH��S*j�lWM?Դ�l�V.���]]]�yyR�I�%3@T��<�P3��c2z�BN>8:*{%�{��8������YU���N�twƞ�u��9j�c�{�t��B�ȑ-\J�1�60��7Ev�O�rgreS�$ޤ�I�"�����SZI���B�U-�ۚW?�ʱk��l��lD_po�� ʹ�q�ܔ�~�J�NCo��8��!x�Z�,Ftϧ��̜��h�w`M�������"�uT��ONmB�����gm�Qx���L�c'�\>����Qt�7�[�\�MH6V^��Y0Cq
���a�/���F�4a���B��6�jX�پWTV��\��4Z/\���p�*�r���sѬ�$�u2>��9_D�mp�M	��P���hgc��QS�u�kӍU�;�
ի)Ra�d��ۮ^8�n����7�b�L
�jL�N��x�Q��{����5��*�>��M�����oEҠ�i�T�%#&V~�T�ږ$O�m��H,��`�z��;ޙ$=�~x��g+���ill4�-2�Wx+���ǲE��~�#m��co�E,���T�jo�v�xa�#WWW�E��;��yX���ԝD��Xo�Ir[w�ղy�g�V-Kjڶ�:�܂�Yy*c�9�T���	G�����gFI��B��+";�I���ݳ����u�I���������|Y����(�ꆎ�Xl��c�gvU����v�90�~�V��5�X]��)f� ����l����pP����rwK�U�,x�J�}Tse)N\�2L�n��7�m�&�z5ZE@6 b �dc:�/d%u��C�,���f �$'s�<O��-x>??�Ƞz1J��"q�L�/
���r�Vl�X�E�zÐ�3����@�1��e�H׶C�
�R�G����]���z��$��rgٱ�n����I��^"���,B������~�R��x�rʲ�'����.���Ѝ�#+����՞,K�A����G
��pԪX�aE����4�mH�w�o�Wݴ"~x�s��Y�Խ3Q�[[�Ve��G2��-^L	��C�i��Th��<ʜ�zl�_��B�[�+�A�������}�i�$���
d�� ���>l>���$��)muj0�lG�������i\
�������%��.�]N�c0��	��S�-(���"������hHj�i�4s��8}Sb�<���R{I�%�&66m�8!Y��������MoJ��a��Y����X�覤�X��n�Cpmu���r�m�]B��=�}.�$�U��!502 a�Z5�R�uf@�L��0*�F�q�����[�$bmqm׬`���ǳlrّWTR�sb&u�,0߀�C�C
�q���}���(��y�G���[حu�X�{3P�qzS��8�O��&$ܰ�Rb��ȗ�p`r��Dȗ!��O�{�#�?[ф��l�ޣ0�s���z:#m����*e��pl�����)ӥ����'f�|BT>�e�7�a}��w�}������ԉ���*�;��N��R rOU7���X�Z�,-�6z����2ބ�-,���̫�jq���7�iR��֦7�����_�D���[3���6���!�73�P02�������|}�u
�!v��c�[1��E����?{2ϻ3S��w~�@�f�8g��*[p
~�?���	�:g�n=����)���xj��,�p� ;�ɳ�����_����MS � -Kq�=7��Ѩ�߫y��vk�
)bl��u��y�����Yh���WL�5]��%"Tp-��7�z���,�m��W��^^�_�	N�PS�*4���U��X��m�FG�95�Ь�̐2�	/
��.0�vZ`le�-�I���y��p\Qυ�2&��0tt�1#1��i�C�(�/��ю�W���J���F�>�"�4�_��L��T����i�f#w�&��ۨ�$[ɪe�;�W�(Skӗ{QP�2�S�?ł��X�]bz�Dn��;�,�L1�~0+��h0��F�/�k��qw�,摫�Jj������P��*���o]F�2�V7ց>3_Nௗ�N��"��g()�*\�>��J�SG0���H�v!I�Eg;�I>DQ�bn�Ji��!Ku���Y�d������j���D�s�@�̡��~Ϝ�/ԭ���B��>��~��U$|�r� f��G6��`����_Z�%9�ے��Z54o�Lc��,��8F����@�ov�kڍ���}�n�7bV�]ˈ��u�I�$�_V.��*�B����/�3��aL�,�c�g�y�[��^U�?��ـ���t����6b�C~Rb\L 2���
��`zc��~p�A>�V��C��W�}1:,M��V���y�=H���B',�Qm&�V�{qWCB9�T�Y3D0����ӈ��ٖ�,�:���S9�hW�J��`�P����;�T�}��6�3<��"���,�s��X����j�*Q$E���6�(�#m��3�f�.>ॅV�>x]�z��>UT�6�c�C��Q�錉"ެ�]�I�CCLVF��"������l|$���C�_W�?dj�.<��t-�:j�g��qde���;�
�ߑRŅ
�h�T 㸓C��ڸ��>�]N5l�S��d�����˲��D�٨[��?H�h�_>���V*H��h��u��p�u9��ˇ:��fT�E����Qh�^�/v���0�H��1��=R&��h̦¨�0���ƿ�0$�/�*�)QUj�}���ivZ$gި�	/��0G9{��3�Ӎ�@�T�Ҕ�������H�F�|g� \��-�kA=xl�kh�<�],�C��6\$O�n��j���!�U� :Z� Nx���ǜ~�Q��^�4GiAJ��h�<��`$����34d��-l@�6~U�+�|�b��Η�7��/s��3�,��;=e��\��@ 0��;���H�8dRh
.��ؚ5�6�Vr�D<�n&E�%OR0E|��o��y(�q�~��d���B�xm��[�,ܤ܎CB"Ȍ��==�����gDo
�"��q��]VqrX�֎y�����Fr�?ڒb�>�[�\��*���WK�~H�Ҙ������^�{�K��px�	��V�5�
�W	CN�YVb���t=S�Ϯ�i�1���F/>�[���	��f/Oh�r��ʈ�������i��oQ�;�x���yi���o��f���L�ypှ�ǊS���[��T���u8���fAp:�����I?vTj5�V���~�T0xM����{�I6TE�me���0v�z#g�I�ʟO�GȻ�R9�Ҭ��Q�Ar��Kť-wF[@��6Q �#CQ�s�"A�a園�ȅ63�z�(�S�u� ��h������7���x#����f�,� p�Ug���7�J+L��TGD7�b˟���N14� �����:�\BQ7���C2��C��c~�����ɯ�V�Z�>�g�X	��A��4J�Am۷����Q���/���A�gӶ �a�On>�A��8������ny�WhT��w8%����IC��D��0�	<��tt�`�<�.���/\WoF���|y̭��t�d��V��]���w!O#<�o�]
4�Iuί��oP&@��l��[|U�=�C�*�z^;�Kժ� �H"m[��l����5����M�o>݇����_��� ����P��c/������Gk�0re&�+?��4�` �զǮ�+��0�ơ������[�Pl�oR�b��i��Y�Z,����Zy��tqE�F2�tvâ ���R!3�@�5^{Vt�4D��^�̭̇s�����6����W�6�k����]c��A��q'F�>��-�K�ul�F��?��C���v�R�J�ίVE�U����Y�/��s�����$@,N����`�O����Ԩ��uG췖Q;�#�SңM
������&��fK��V�=��u���`&;����/��~zSV=%ʊ�=���'E~;���͚(�e��b��~���ћ<�<��Ej����йj�c۲��ݡ/;�g`�����6��ӧ�i�h
�<^pe���$!7�`�ē'��\[3�4����5ۦ�7������[�k]gIL���l��K�v͂O�C#���!^�BN��pAB��s.���ky��y�Jf��������.Eƍ�%'�m�$���7f�}7��^�w((>O>�-�!��Wa�L6"�(���f����%i�D�$W���K��Č�z��L礊�КW�Eˣz��x�P�\%���·}᭝�8%L����~L�6����u�{=�XE���NiႏJJJ; ���7��'�����-d��x�����?��۝K�����]{>TP=oܤ��Qx����q��a�<���|[��?�ӵ��?b93Zx��T�I]��b���뺊�oaL���#2�q�E�ޅP���Ý6-26o�bF
�}�:/&C��\}Uz��3n�P܄�7)�Zt�u�e���Ĩ��]Hw�P��r�����;N'm{�g�2�/�k�Z����L�(<O��(�8�׎�mOX˭���ej3j��]��:r�.������?82X0�^Q��د%���Q+����G���x����c������탊CכUO��Ӯ�gU _i��WV>�F��l��N#V��#�W#��3��X��y*�U�KWi�7�JX����V.��\�j�bj�I��ˑww�PR,���
 ��o�|�w���\�\�E���x#F��q����<g͕��;X�`uQ��^��T��������g�C���nTO3TO��-L7�K߆^q�u����k�����z�G�n???�Ӎ^u::��aн��g�	ɎN^t�>�k�a�҂���'���U����cS#%" ٥/��*�$x�/���2�T=�۪:҉�����L�����zv,؇��:�nV����_�c�����atA�YKF2�4^l���!xN����RK�� ��V��gHA���Z��)�9�^� w�1�\�ы��[;:b�8TTV6��!���*'��eu=��h��ei�?=�1�8�K�������s&���AY�҂���F�N�� �����k_�K�]���˭�{޲�L��c¡�=��	Dzy��b̖-#�RJ0�j��z�:L՚���]:�Z��>�8����0�~�ˍZAp���kIL��D��j4������9V~��/��NWEEE��t���ԩ)ڴ�h��Ԉt�+~�=9y�ofVV��/�a�$��pIf�)�	KNA�ؽ�@�֧��u�����#~�^obC�s����U~���2O:���f�����W����w������[�˭"S{;�'��z2K\�I�z�u�ф�p��I7Fmn�x���_�U��~(����ϕ��*��U;�*�B'��i�i�E�K˱5~�ZD ��(��?�U%W�T��_������d ��gj�P�!N�D0
��&���`!|Qͯ��a���
�k7��'�"�1��!H�2��殓c0��>Iv�]��+Č]Xk]*��ciɇ��h�  0�g~�� ����J���{E�lf@�4�"���� I��4Y��=�V�F}������>5�Р=F��k�P���	Qj�ZC����� u�m:�����4��������˔&�D�q�s����G�{];	,�q��:����Q��C�Z�s��狗�&����h����CF�+���xO�l'��;MN�l��jq��<�W�!��H�Kf��ݥZ&���0qpƧ���S����a�m�;?J :��n9�p!���dj���/K7.�**O�����"F^���%95%�>�ET�t�.|@��v0���F;\�w��P"��tn�v���"Ly���s���.��%���^r�伐D;���5j.~�9���Ͻ�~�j�Ȗ�e��J� ��J�e\D*&��Q�d��-�c�о��B�� ZQ�K�I���
�4�e)�466=����
���� �+��Eժ7�1m����8��j���Pt�= ��>�`�r��e�bgʵ�kO�9�|�_�T+��&D�͟��Ω�[p�W�E,�<�K�37W��8��)ˑ�L#���lK��7�-��h���_�~~��GIôU�L�e�:�>��b��E���6@��=^�dN{]�0��O)?��'��c?�Н ��Iy}��� Иf�D��ԉCDE�7����
%pv��P]�/�X�4=^���?���K���4,�����]2T������TH�y5~���F��B��Ae�O��w+åMX��/���"48�$�E���*V|�F�'#̮Z&z������i�Q�\o5��<(x���.[{�2#��;kb� ��������!�~w��.� ##����>��%
����o)�Aw��)sx�_BL�edZp���>X�K�Z�a�Ί��G��F*))�n0}�f0�#S���fp)����^^��g^���O�?���>����_�7у�dʝ�Gqu���B��G����c�P��d>䄃ůt��Z��)*��n7#�Շ���Ǉ^L�P��/� �k���p3u�3�eK��%T���P&��ju���"�n"}��Z��J�m�IwxG�?����`�jܸ�-���pՀH0�2o�Y J�+ꏟ�S7�����U��ߥ��2}pX����Ϳg�D�N�og�t��3-�0�&�
��7��՚�&<Q������b7���E��>>�/C�	 "Q�	0A� ���������>n���y��v�s�*��QX�\��c�3��w�H6Ġa�병���=�I�����S��@_�<�|�a��D�(_f�I:�!�&���*�d(���ʞ�e���fA� �&��|��Ȳ~������a��/�% ��?>~�[��h�Ώ�Q�FYz<���F1H�؅���������9˥s�9њ>�w���8Z�Y��ϔ��i�(Z7�y�˔1>�w!#�ϛښYFyZ2��� ɔq��}^�8�JR�J�j�u�˺�d5����2]pNc��A�0�����5���>���~q�|�Z�DlJ��͛����\��_M>y�v�x�|e��-5Q��F�wA 8e���F��d��r�?�0[�3 �7/7w��s�Ոs/_�쇜�Cv��Y(b��L�}�l�+H��?F��l��G<�!��ɔ����!����N�.U�xΫ?"ՠ=�W�u9�Z���G�n:y���J�Mf���+��R�"J���(k|�|�Ǎ`$�[���ܴ&���P��sr��5�̽�����6�-q������X˾w������.��:��<TW��r���/w
��}�c9�跩�?�=�4kT/[C�:-N9�Mb�^�:����NS=�̦r2�8�ߴ<\&�a]�~+3?��;.��յp���l�ۨ��G+//'�p�n��U�DG�ǡ�fl?��
 2@t;<�/O?���ގ��/�]/�~�^<��+�*no�=��X���:�ẵ(J1�r�}�-�H<�?₷��WC�ڤ�\ ��ۘ9@.��			ٯ��M��((�s��t�����(sd������ʴ��}�E?� �W[gl7G/��qD���i�f;?Ty�P=V`�PL,,S[�(sD���}�Jo<���$ߞd�a���!�_󾢒��[�+�p'�*|(���ů6��랯�8��y�O����V�6�g����zo��aK�pU�;Ez<@��^FB�^X�������T�u �����~�W��_��R��L�i����L'��'�"����8���It-���$����\^_�Q.m�0&�:�ڢ��l6�w�LoNV�fs��"p����	�y?��|��t>�tDĵy#�� TTF�C�~�=.�X�I������d��k����3 �;�����k��̾�0�y�ҧ��7�ԗ� ������/�;��r�F�Ɂ�f<E=�C<NV��>���[?��AH��ܦ��_T#Yb���q@]	#gq���OC���0�Mg0}.���a����h�L�M�j�]�0�K7g�o��h����;���r�tI���z��[α��q�&�X��2���7���rs�yZ������(����d^���m<��e�V������c4k41��!\o�1c�W�j�m"G��0�g�7��Չ6�9\�m��-��M��Ι��q��Wˁ�4E��hd�	Sa4h|盝��J�a���|�JJ}5?l��5u�����IN�`H�����v���g��1�}l�>g�/�R�K�$V��<���,�VVE���`����ó��G� �O���N�?�N���� �)%�U�m�\�dϟ���q��N�ct����.ׇ��1)py<��l}���ە9��F(����� ���tx/�G]�謍�(V7r��Ϧ��q�u�|͎�{gs��&K�?�1"+�d-}M�f� ��I���J���Z6&}r��y���;Uzϑn�h �����Z��1fc�� t��&!��F�R5FF���9r���H �K$���E�KZ�By=�m>A�[_�MWf#���4�`�����ZZ�-�!�rDZ�᠋���_��n��O,�w�#Fi���Y�G~FٸG�Z��Α�U{�*QW��s����|��0!u|:���9k�O�λ�k>;�8H���C��"���X�ɠr���@��G��UF��H�w�<~����-�{ ?�A�ժ�|�������BD��Ԁ��&��~���G%w�dɮ����tM�^1B�jmz���}�"C���B4^�\KyLIU�$b�͏-Y��?n��DP� �$b�ڢ?���V}�G�"�0Ԙ��i�5�l%-H[y�\�l�+�_/�~q�8nf����;�;"[󳰷������ǂ�+�7���O��S��X EJ7hz�<������	�y��tx�*S�" �*�����|�����N����#��m����a�߆ B�9M�{]�O��s��Ȱ1@�y)�k'�s`� �"ʎ"�9@�R `�h9Ef)��h4�5󶀚qui������0����7'C���l�7/�.%8
w�AV0�>���� {F5�Me�`^���q�$n^��_$3w��^_�|���ֽ�V{0h:��k��׆� G��ȿD�/�]��?���n|'##s��rS ��Un_BG'3���٢�ע���ӻu څ>���ހ�C�fcL` T��L?��ձ�Eő֖ cU���IL��4��m��T	�����4�&��� �VΥ'�����!�R�a�����7���FY�g�7nI��s��ŭu�:��s�Y�,���}�'.4��Q�v4ub��<�`��1�dT;QP-�a�{���i6����Bo*���]�~1F����ޣ�^�Q����|������ӎ���G�U�w�K:�����>�/���EccQ8B��[������r���oxS^��hu�3/77�,�O��J���<d�s�XNo�T�e@U�)��]�h2�t|7
�� "��:�[q��{��b�JU�J��AW�rS�3n%�x%�-�If�В���տ��S�N]���������<H��a"3OLP �mD �Y��9�D|/#-]��"FQ}�T����8���c��^]K��T�t��B�3�Ԫa��V��2OW>O�2���f��ټ?��bܧN|^������V��Ǐ8��	�����>��۝���Y�W�����}����nX����|<xuছ�1K��������O	���t������(�"S(�����QL{�y�L���#�T��ҿ��c<�9U��y�ϱ����re��ds]�P����S�Y��6�m�C���D[�W����u��4�k��i�8i����аg�&�[.B!n�A6�������v0��P��z��^�;�̞��m�]^]� ^�&�ǁ�8���t�qkz�-y6Df#|_��n�;K1�E��&o��WI� �1��dJ��>|-�ENɐc���Q����u���}�iDV��I���礭�;Q%V���x���I����Vv�������c"��2��o��x0{�6^��[�F�7�Bar�T��U����O�AȰO��������~d�b�--����R �Ah�I��@f���z5$b���r��,���E��(�3�HqpcEj"�oxg�T�y�$���UUo���T'��ɳ�PM��j3��d[;�T-�a!S�1�0R=t�"��$j�,��
�ɦf�"Z���\K�@I,��o����[B��%�B23�q�7|��+��������v{e�Є���N��w�h�2<i�e���>�U2��� Deա���s�z-M�g̙#�+~���#�z�1��ԋ������[���B���h���?�U�!�˲)I>�3W!l�pϓ�(5�v,V[�nQk+�o�����Q���>���,"qvd|r��1+R7���W�X3G��X����;���q>5�\Jm5H�R5;�D14&���P�|Z�����&�0�&�v;l�N5(>"`9�`�I��.�NƂ>`�&?��l�7��)a������61�F�ڐ��0��0���-�ii��pr����D�u�	_�泌�3ۘ��z�����
�Dg�5g2�~Go8����&F/��"�����!������#f����OML�],z��/���$(&�CaȂ�*	n����>t�ja��M�Q�e6@-i����`L��|3����y���q�m�8�4H�)c��!j8�F�<m��7�@%7��H�-�`���5ͼm4WH*M:q���!����֕�SH\ƞ8�L�t�7_=8j$����nK�$�0s���,�~;_ޯ�Z�5L  ���;sWmN�?��1x!��>p�H��͟�V3�!$�N��t�]nCk)eh8gnm�z ����l�yҩ{E���@�wb.�8Z�fM�3'�K'���=l�Lߑ��JY��[ϐ��5���*���/�
j��Z^�X�əS���7K� Bl���IDѻ�u�n��
��K�!fg�����?���RM��I����1�e�v��X���ɻ�r=���on�g��渣i�mpX��'̫�"�b!!���RE��o��Y�9�G���U��/c��eo��H�:'���%:�'e9O�!I�����Њ���ѱ �M���'7��h������哎�!AWL�sȴA�T=!��n����!�,�Ud�{%	#��Tz)	)7�h�$�mo�5�f])ႌk*M�_Ҵ�e��e��n\�K,��|I�1C�^�5�y��
�����_�G�uW�+��<�Y[{�.on>!��s>>�ɠV�tQ��g��~�wR�B��*F�?I&�A��6]��F�JC��c��fq�����H���n����r*򫟄ﴠ }��{��}��%z�O�Bߊ���9��7�r�����"���@�#��#+U��)X������G~tB��۾��813}-�D�,����7A��N����U�'}癧�ǽsu��)a?� �������ǽ��^^�����윜�:vcҧ�'U��/���^�ٸ6�#��Zr.ߜ�H�sTBp��f�l� l���+ר��S#���k���:���2���,<_��{X&Ơ᏾�R�$�8�$5&a2Uz[�n!Ǡ�����j^��)� �C�>k�
%�ݾ��Rå�t3H�7F��k��c�íz�^�k�ۏ�Ŝ����m��&�u=ࡾ���T���'B���9��`��VB�7���+ˉU�6@�Q� ���=���7��
o3�Z������n�����X,~\p?hd�rP!1����,�\��eސ�pQn�5%�Wi��4����s�X摨v�_Ւ3iZ*�se��������Z})�~���қ�����S��k�}	b�an�P`���X���rt:�ep	{Yr��X��ͼ�&#��mw����O�f���F�აG�g1p/��,�?~��0?z�Ҍ�\Y�ci��K%c^Ҝ����F�tUNx)�����
*�dz�m��C]�d�ō�Bh�z����`]x�<��������	-�p������m��H}�3D'��X	+}i��d؇K�zɉ���὞I����`��n}��x�۹
���o�u�B�5�~��نb���tI����霻@� Dd�i2��/l�*��L��
Ƣ;aC`0�q�Wa~�j���7X))E�����W��BٿN�Ԙ����XJ�A��ÊjF��{�\�y:h�_��%I������e' S�Kp�6�&{���0���	��SZ8��/PJߕ^��\5�[ڸ@)�>�$K��o��~��(�=4�͢�wYρ�U\ErU-�1-;C�=0j?On��7���c��;���}�ҶY��BAЗy�䆄�����A�]��r���Gf���!��*�Ջ�\���(�.6������Z����[okD7rK4�����WK�AX,O�&��K� �*V��ldO(}�ER����0��½�{Щ���Y+�&z��Un�te�Z;�C����U����PeK�{5�čZЊK�+���܄���y�/Ʒ�,
�
D���C2S�02XHc���R��u��9o�E��:n�k�v_R�h��J䲃5T�3�V'�ͼ����$�ʎ�Yq�>B����A��_SF�)�rV,llӧ�������Q_1H��U4i+���nlҧ��;�#��c��c�
�J�$��^����hE�N�Guh��H����1J1(����u�3{7���WN�;��߄4�0(������vT;^��O"%V�׵�U�SG���tդr]��2W��{gV�;��g��n��*�%��A',P�r�	W|�����&3:]'u�� S��&�=��fz	��6Gon���D�U��:~�t1X8==}�l\:�w�Pl���A���b�	��V��٪�:ez���e�|`v���.�d��%+b�<l�|V�'�廬��d(�9,����v,�s�(�fm�=�Z����O�,=��i"�$��@*Q\'����PI���gMwU����239���O]	�o����U�m��kmU(��ʗ�#�l��$/�{��(�r##R��!���рo���E���K0X$GőѦ1��j��mɔ'��i8�~�����v��� <v}s�P%+�����d�Z�,l���]�Hi��������k��������Fb7�%���[�O�#�Js��*��:�l��b�4�n�eݔ�&)�h�s=/Վk�,�l�r�W<���+u�\%7oh{����L|����UJ�2���9�t��%�������\X�d��V�'ޓ���8�}��섯䋘���D����j�pO�<"��'�_b�� >y�����P��g�s����Ƌz���&�1�\j/Vl}6�|��� �*OdU�K�����^�һ9�^�����L������k���I�2��N�Xb`cJ��W�\�C��SR)��<�:w����M�61��4o��Gއ��p�(������}`7�����qM��r���o	+���U��;\ҟ��׺|\v�S�߬8߬V(�����r"���֒+�'RHx���)�U�	��=����E��l(�I�/��94��Ȑ�NPks]��rdlgg�t�|3�[tR�M�"G��Y��5+5�w��y��_|��,+��h�v3'�&{�]�8��^`��6f7���S��T�f�Iv|�"0?D�B��f��K�\_�DS��,H�U��W�=N�lڅ�>����~��YA>�O8A��z�XA��vC�#���{�*2p�p#C�Ed���������w b�XæF�����ʍ5�B���P�{(�	�K.�#�nX�;��$=�W5���iF�>h�O��	\�(_�nB��[u�c G����iT�*�����?��2����-��;w� E�;�����nŋ;www�Sܽ�w��3�L�%3���9��n6~6F��6�5�͐R��~o�'ǗZxh�,0`��������>�?tl����I�{�v'z^i��-�~*�����5}cegj��w�t��?*���1A�Ű�83�m�'w��I#�ad1a�ы5��5~w��]�߽�a�6I>�s%铃Д$���3�~����2�.Ȭ�jɤ2�;��$�I�6��DA>n>;���Ӵ��vˆ�wIq�����Z�C�>����j�N�����AT�̼��*<�0�`.���6���;>$��q��_P�9�Ȣm��ͭ�7n����\���ש��5��w�+ɚ�	DM��-�i%f�Xq4�W�_>q��%H�������N�6��0z ٯz��|�0]�CȘ~��۞?��c���� �+��)N��'����qY?���s�̲��|8�
��O���F��m���/�������n�N8��P���3�~�nFh2�v2�ʂ/����N�D�+&^��R�|ݖ	<��T�+�n&)�j��:�EM�<ƱH�<�����Z��c�k���T?׭��MX���i��̭g��-���bVLL̝���V�EyE5��G�V[�Θ����eG�mI?7�<p��m/�я?��8���� �>�L� g>�~V�?�����j,0�$Q���b��ᮊ&D�2�ڏ�ܷ|�YZ/ ]���?}���b#�{h��ˑ���N���������"�+�l��?��T"�y(��O\,f1����̈́�:���
aɗ�'�O�Y9-i�fѦ��&K���DCz���"fU�:��f��ܞ�����K;F�ьZ�L�Ҝ�բ�G����@�Yw�s�>�jJ�}+g�[�	����$��B1�|��$�5��7Ǝ|u:�]�j1f�j����y���.m2�)�>Q~�"F�%ݎ�p���OO���͕�lB'&<Tht�^4�oZ�B�_N���M_~r^^$Y(�t�tQ-4��#�<��`���^]N 5�5�}(}�I�E�ՂAt�JN��׊bZ�'v���*4��C����4}
>�xTU`���*��ւQ�PZ�k�V�S[�l�?X͈w���c�����;���10,=�N�2%_�#CYUʘ
�2(��<T���g6��c�R���M�s�0���w����ZUa��if�{�ggg�1x(��6��!I���E��Lģ&'�{Wxudk�UkU�޺��̒W��n��n|5��[6C�zTkc�\����݊m:�:�1w�%��ׄ�p�k)�J-�:��9��m�V��(�֢�'�8�?먛
"��������^��]��=��������ml�'5c-/Ӫk~wI���ԇ%��ƨ(q�'�ᱹ�=��l��O��'�H]HG���o}��V�T���M�.��p+�M}�n�A����W27*���5Uh�X�I/�Wi��=B���B����+d��2F}ʍ�O� .ҬA�f�[T|�]N��ML͋X����+����>����<�t���;�'VzOnK"�q 7�@��(�]��i�A�Π������'K���AN5I�;)�^�7�7���0'W�L����pI�6zO�	} Շ�I�VE}��T�q��w�{�e9)LwA�`u�L�P����б5�1͟H�/������32A)��d_��CW�dd/�OK��-QW���Yq�7O4K�?'�۾���wA�W��L#.����� !�^y����Q�쇸�Z���f�g>Z	�r�(åD�*m��m�Vz@H��a�&Ufj�gc�$�?�c3l7���E�mPK����pޱ10JH��Q���R�C��sΡI/4v�U�Y�@8��z�Ψ�����>v�GD7�9�S�b�V�3����EDt�e�+$��BA6����WJfPw�ŝ�q�79pT� �d�^��V���̖76����Γ��D��H� <axs���""��.h4�M�`� T����ϻV<���4y�YN���t�׋bOJq ��+�p�~M�*V����+�^ӺG#|�uP�ZVVó�70�G��㐦LPvXe!=$��xq/�z)a]=����m��EI?x	��RC�F��C�E؜m������ؼG)x'�v[���$������ɵ���TʘiJ��X��+��d/�l6�t�Ro���ΜWD�T� ��T_;,Bn���v���G��fȍiƮ	����q��b�o(�ڌD�'�v�1�&�8]~UY'sr*�V�ԺU,�wsO�����s+��G����F���֡K#+g= ��8g���X.�/͔0X���v�~%)J���b	�YH�S�D��B�	��L~�V�<�b��0ɟ����]�.L~�A����*R��#�Bq�Ԁ�к�3&�b�P�Ee�0r_�y���������o�"U�j��'#�YF�K:S��:E5�1$��e5����4���͌Q��,��9�����5�&�9��ť���w�	ܖ��D�S|`�[�i�^`���{��ʋ�ZY�բ�"�s~��s�A5��By�ߗ����[2lȠ�MI�K>��9���<���X�D��U|�����J�ƿf����&��*Z.��?W�4�T�!�PEz��n|���ŐG|Vy�@�&}M\	����W�K]	ھ��Y��!��0Ox)����S�d�r��/�KKO�4ag��8FAH�\�I��>=hsu�PK�������|��e�S@��Z����;[%�}�U	ބ<	Jn��0��B	����f�n&�;�vd&FT1oE�e������_i�*���l�-�����l�=�[��ַ���Da3�mfw[�hu��"e@�V�ş������P$��M����ҽ�M)t��ɳ��Q��S���) �h�j?s���ױa�Cx�+�bb�Pv�!2�o��b�4�;SH��(��\ ������W+������8���885�������)/�v�x�����PpcH�1*q�M�Q�*C��JV���1�A�2j ����碉�o�仼5hd+��k豟sc-e�[����~~A�<�Ċ��:]��8��e�%:s�4����+������6d�e�f>E��u��[qk);�pm��x�6
x>-g�4{z�4"�s	���|��(��
a|�f��H0�W�����{�,�� �x;:�ggg)W�����LOO�	��e�r�ГJ~>~I����,�锚�Q(2@��s�"�V�6��z�%[<��9��>N��P�RZrRX���
�L�7���2Lǻ�d�|�*\�?nOY�a�I}ϑ	*K�k��V��ϔ�+�a@(�pY �`�M�d�CN������Y��XY?�s!�߲�2N	SX<��"e\hJ�������b�֨�}�����sX(%c*i�����L�M�i4 IСHOɫ/LL�>@.c��D��!ڸow��e̬&��L����-�ǅ�H��}�e�m�͌#8�?��d���H G��
���	z+$߳�zy�#6K�=���3�v��$vvv��sGYk�����ٞO�4o(Ұi�g;����p�:�l-U�Jb�^����"�(�siBq�%�<
^�n��r�l�N�Z�$�e��t����j���<ȅ�-����.���,�!:\���9����(�o�p���*����ꗚ3����\�$s�/Nu]��d��\/!n��o�/	KW�i@2e��)�x��EmG�x�h8�X/Rh����I̤D��u ~+�O�H��0��t�/��W�4aQk�O����H�5��]��β̠x��3�!�����@�U��^
���Z&��f��I����0_#P���������	tOM繲�~VF�/��H���Ł��V1�T㇅�D�e�>�V��-JԚ���z���T�k֮�8]��͑}e0XS��F�����س��\6�~�Mx�Z%ڤU�N����6ď��T�ē���Rݼ~�q2�C#�:SDh$���l��A���[��ݩ����`�r��3rӠfD:Rq��.8`!�g�r�r5�=&�U�[$c,x��},���L���\�AA$�^�Y�뗑�\�kĊ�?��O��?�vGHfu���<�z�Y�w�>�������D!{w"��3��]�#U��`� c5~�ȁ-d1���܄4�������k���4�{��5�{xn�Fi}KW�G�.�LB�|����O�����>e�	{��MQ�Φ�ҩ����ܘ���'�Ёr����������}K�䜢Ф�_���ЎL�4�hw�`T��S����8FZ4>&^�ɹ�*Q����{8����v��*�*y5
9PX��I�,���L.�]��A�'A�\��B�g|c�0^%s�����S;��F��K���e�"�\�+�D>�Y�&�1؎��ʇ�Wڗ�?��ie��>�M%y���	�������Oeu���h�6��-�X����&ֽ3��|�>��# -��ypԈ��d�������8^��/��駬� bTC5d,���V*؉��{vYr�!T���P��J��x��=�0��Q��h-����R���`ٕ��p��e��'��m�W�=龍|n!a�����wf�N��FyQ�����B�H����#����X�v;��4rL�s���N"�q#4=S ��zj�"WO���ki���3�M?����ܝ��aM��>
'��D�ј���a������X��?�ʒO��Z2��<�D��FiմRs��O��Ef���,�OQ����>�BSE��ס:r�pd*.&p�̲%X0��΅�Ӊ�T��6>��gH�J��y�'����Yb��R�%|������!�;Ӯ�юfûg��%J�H|[�G-"Aِ�0>T0%����Ȱ����8����CAD���w8Oն��=&F�U-�����τ	�?�K��UW�i�>Bg_ۨo�k�a�
qy�;�	b˷���ST��"�fĕ��r-��vN;c�_r�{yB�.�.h����q���d�k+#��R"~9Jǰ;Z58�
���Y����f��ڀ>��&�M������|����,�c���a�9�nWE2��K���$�K�����e)�;���TF���,E��7�v�h	����{q�E���nإv٥�9HUC�vQav~�o��o���5K7�*^����!�W=�����4��#�Z�'���|�(�e�3�,X�5�&��9��p�X�G�;o`��6'�^�O�6if,��4ØOe��i��!|P��s�V?+��
7���B[�v�W��i���<�T�@����>��:!PF��=��i�k�2w��R^����V!���O�VY�s�������.�PL�gEs�h�tw^��ٶg@|ˌN�(��K����dϋ��ǁ���%�W�t������:�._��(Fqs}?w�[g�^H&f�O�[����5��%���%
���ar
�Ŭ ���g�V�3���R��"ٱqp4S �7X"�f鷯��w[��U��|8?A�[������.G]h9��E��7���c��{��^� �X�0 'Q��$���rk��[X$ٿ.�qvx(!�V�~g A]mm�����F����}�m�(C��Ԅ�ѣR�N�X�Nk�C��uB����P��p*���X�@��R��g��"[�-�����>f�B�g3i�-lUKxal�.歝�T����@�7��z��;_�I��Gq�X��S�e,��۷h�^'���,,��#ۦ,VE�_���x�ͮ�F�Bi�������
�'	� %{6�g3�%f'�;�����k�XkC�1T��O T����{==$�%a��F�_�z��]�j��LԦ3Y�	�I�%ʖM�|����޿��W�8���Ic��-K���V��Ϲ����7d4�Q?��fg����z��B�I1p>@���l��r����̖h�����˶��2��3!������w���_�η7�H��kM%�6t	��@"�W��M��Ժ�ʖ����K�n�����
���t�,	�\-}�?��sICW��}��(3�sYo��:����&
�Y5Z)�a1q5��*g�J�,)ٮ㻳dHZYx:��U��xC<Os\�Nv�/[m;P=7|=�����e���w�/�~~9�~3`5psK�����Tf��v"�쩾��!O"��2k��]��(о`��N@�b���������y�#�^���NJc�ؘX��cƒ��R��Kn�9�HhP{{{S���^A���u4��6�W����E��5,]�m��|㾤��dV?+�-��.��/Hz4AJj8�Aᡮ�I�ӯj�P������`]~'��͊d˫����s���֯�,oŖ������I*w���jc(�YߝÜ���j�}jʭ������:`��n^��oR-#�ҁ)h��j=W蹴ç�C��κ�ԇS������<��X;<,:_�c��M��څ����\VT�U�ަ*Td���fU����Rs���.��^z#�2���I7�,�Fs���0�ѩ�u&x��e���@�7=��K�\���PD\M�QYW�މ	9A��/��q=�����|����@�a�06>>�O��	��L	6��5�ft<i4�%+�t�WZJar�D����/�.�Ӏ]��a�x,��R�KR1������dvD9��{�{�b7PK|ފS���<*�&��?%}�+�nys%�2�,�(�a,z .��[���.���-q�T��8�����쁍(�U��#�Dt4���/��-V�6�-�Sf� �R�ת�(�h��yY	I�C̯d͖l[�wߐ�}U@+X ��h	FDF��{7�ws���+���鬝���[o�����?Bg����CG�|kɽgXU�٧o�V��˒���j�����2q�c�.��ոȞ�ē6�~L82 �=������,,�{�C��mr��F)Q�=8i:���@�i�`��N�[��^qBdPN�9�b��Қ��_��.o����<�
s`��t���ʕ�FZ��QY��!��y\m�;Q�!:Ȥ�Z:v����<Wb����~��笋�=n�)2�)����xl<_E��K]tj��YA�H(�V���G)�,�LQA`ˇ��R��í.Ǿ.��*$�]O��0\��*6��ۨ���*{��yif��_�F��Z?�=����B�����)�Ｒ�F��"�h�{D� >�C&�r�]�����%,'�P��f��� VnS+:Ş=ňˬ�}t5�YP������������e�<^���#�h�����+��d�?��M2EF�I��s��C~|�zD�e�"���L���wN��&@f�m`MnLf.7�W,�o���Վ���������F��~b��)%t�*l��'��U�0����0�Vt[���ew1����%J���M�0:]�}g����7Eab��hƙ�J4sN�QL:S��ʔ���}�����;���F����r�'�~g,:�5����"�V�1I�q��)�kң��Hǈ�@,����T�9���I��e2������rǽJf�X{Y� �h|'Y<`z&	EB���.ϿE#<��y{G`��M;�e�����}u$=����^�ނ�����Hk�/Ɖ��Y��f\(-�)�HB��hvw_��عU���<�ؤV ttps�n����z��s�8���ƭ�D�l���nuuӫ��'+U�C��V�D�ПN$UjQ�77��|[Q��l���2�y/3�8{�zz�¢^�g�j��a>����4��F4- ��W�6iU]�E�Zw�6���i�A�<��KI�ڰ7`.�PE�Y*jiI4����� R�A����sv8��w��$����pc���NoY����%�)�w@��Cȳ*��S��;��4�9*٦�w���a�� �296���l�����/���g�E4<(C����}^�V>����M?H$��/���]�gx��zV�z{�np��[N,��-ZNMV����L/���2{��X�����o����z�ۚZ��/9���W琧�X����sE3Je��$Hr��:2j��Va� Vt���z�'-6�R�F}� `S~� W�5�0������c�g��s���r�~tq�F���8��X�e�>���b5���]�PNY�I����F��NO����|�����#����X��`G�����p|z��g�P��O��K��,�,��+�~8�����+��ΝoW��.�x��JԮ����$rp$R�ZU��:QCO���&3�8O�b���*��m2��<qpy]��,��!�l˙�LCC����t	�%�����Vy�ݟ弌LL���?��G��	��wh<��G�qYu�!1�"K�7 �7����9(η�,*Q ܰR8c�f�l�
��_����8A�v�,Vtl�Ř��d�a��Y�o)Ɖ#Io������ 
�zd�oT@Ѯ�@֛T��ʜ!R�>V[�q28c���}�T��@��'�?�j�ff�H��K�^��'Uj�4�UUeLȎc8���t��~�3�h��'����B���0���g'i�R�oJiӌ͔T�T�	�X��(ƕ����Y��6-G��*2���-�h;2�#����.��&!�2�^\���=��{�����j�	3�HSn���<7�%�:�uZ��ύ�P��B{oDC�Y[Z�:8�vZ'\yU�9	&��de�� ������ʜ�Vd�`F�ci,#M�(-e×�#l3Ŕ~l�I�&���G�}G�gJ3�˭�Xg��]=d�v�ғ�e�T��tT�!�ML+3�B�"�`F��v�Uwqi�fz;Fo�*3;[\fԄ���-vEq����-ަE4w�_;��L�� �sbr�HVx�io%q&d��By���a 7��|`4�A�VO� =;�<U]7ܯG�]�SjkcC���T�b6�b���E �v�-�;ᚺ����,����($��-��,=��
����-k��,]�CQ��Mkm~5⢴��*�����p�i�A�s%�q �����$����;R�i��E�Y�VS$x60)n���d�`�;��{s}��{?=*��b
]>|$�8m���l/��-}��x��W��wl�/..��Y���D��#�U=�gi��Y�`��,��}��o�xa������`#G����:\��gd)�*���.��*.I5PG���7s�GV��G����� }!�)uL�����;�U����H����X}���Ł��=^����Bne����������9�u�uLB:6�ē��
�B�[���&|6���Z�6׈��R�P]��w�֩�]�%9O��~���4�g�j��®%����BSs( �~�*+x�Wed��s�֕�!�5�	@+W�t#D��?�͇n�=�{]!�����ߥ�B��B7�/B�Q�B6���'Ζ��x�d��H͖�ײ� �8U<Z*k�p�z�_ �.�Įl�|R���7X��m.w�4��8L�m�����nt��ݑ�ib�AIA�%
{qa�jjjx(�|nѩ�O0)�u���1�@�ؽÛ�
ܧ�D�@��P�?��|0m~P�y��;>;���H�4�����>DQ��޶>�I޷�^�1����]�r�������_��ƀOT�n�f� �*P�"��Xm��a��PQ|FڐrnW�����͋ڏW��#��읺Op�������_+���{�k;E�)�N�s�<��f��"�<&�sd�,Hk�<vO/T��$�(�򠜞�����y��2H�ea40�]7��	�r�)"�����"C����?̐�oI"��H��X����N�kQ����,o||\�B�\s��O{�Mv���u���4<�����GՂI��������K��Q8��[z ����B� ��7��׷-����s[�ic33j�20�8�w�w��Xq{��L��<c`pޒ�3�1�0@>��{��=W�����0ͦ/���߶.������o��E���z���<S�,�h9�8n�n�n2��c�O�+q�[��R�Z�B�S�9�BQ�v���T��e�.Ԝ�?O��z�#��F�^7�u`k���Z���U7����j�����,�!=;{�N��gz�nGeކ]}#`��:5b�Hljkc������5��|j���z��cy��(<ׯͽ*�������_��`����z�G����.�F����șs'��'Z�n�KͰcE�'H�W7tv��>��x]�0#��*~L(*P'�O}����v�%��Cb�����1v���`���j�+#��Q�~��&<�t��*�G�V�� S������Bܦt���Y�܃P��,Y�My��@��ŭL��@`���9��fۃ���^X?1� M���	�b�aqc92�߿��O�o`��QcCO��0���>�����-����R��h���������'&��>����\*��B������ǲ�o�o�F�����H�1=��MG���Y����A^]�{t�c���7���S�䊝������/��ۜ���Z�W�y��w��E�N���x�e�ic!EG�!����vz���/�Hk�AW�m�=E"\�P�����q�D��]�������?=�_/�\��a#|8V{]�ߧ�/����)�z�%��F��v��E�g���9sq'�縹�o���_�������9uey���9�2���qin:W���0�I���ˈ�ʩ! ZX�g�_����pY�� `bݪ���n�����}k�S4�8��5�6�C�X�ؼ�t�� ȐT��:���{�9#��T�9����Y�(5�)�]T�$��	����a������9XǨf��/o��'�����p�����)��"�����ҳ��xM�K8;?G"��!����Ifq�9��B"(�4�����WbD(z��P�`����%L��m�l��P�Y�S����f���`��[!o����$�{.@髻���`=;��� �VEk��vF�Ix�u�(����\[䌅X�M$y�N�u��S����z��嗶3/<��eHbX�\��U}�;]����Vw���Q9�454L|}���S)c�&��[���m2����;�ӛ��j�ܭ.�|:=�17�Ij)+]�X��y2������:f�-�F�.�5Tl�$�/� d#�aT��a���n��>��Q<z��"��S����KTD1����x;p��q�X���`�}�Ǯd��1F��/����3
!#I �/s�X?:��K��l�"����]�|��n_����+ǭ�B���d*"�]u:
�ֶ{q����4�����,�9�u�XŇ�II'��D�K����	����=�u^M;�g�\ߒ�r����=N�N;�7�;��V�^ɲ��J{J����`��'�||GǙ�j���J]�l|V�bKQb�r����`A/oI/��u��9Wh\�}�cĠ4)�j��C8W�Fo,-l����^}����u������y6�\�ް;�_p'2W��o���R��3��F�2���S�Ý.���l`j�u��O�����a��N�9�����?�P�P�6�0l�1���1X��>�?0k��2Ŗ-��,e���0U�U�hi�n=]�ۤ8�ʚIcK�֖�A�p/w�J�A��y�m��c�>���@�$׾Lābɿ��;�*�*���HH���_�/�jz�s���{�6/p�}�5����GkÍ3���t�N��F{��>Htۜ��@q/�������[�^?���<]��vݠ�c67cYO�F�T�z�-�0�L��%��:CP?�r����,��U5�������sm�s�"���B�����@>c��v0l<�H�,�nU%�Q�m�CXN;Tf"/���a��U�2�(�KFU�]C�bL��v%0L�i�|�+�
m6<^�]��4=g��u�j�D�����7���*hOM�\���-IlͲn`g8���r��p�@(�8��s����<�*[>��/,�S��䘅�{�����=�E�=-	x�}�������(�,�U	�by�g�%�b憡��Щ��
$]�1Ԡ�����rI^�@BO���#,�o�qY_ �:��]1�%���}��V]���/��1h�D�h ���92\�g\#����ttb�"Uす�gUL2S�>�`���44*�>�k>hˀ@�_*�3˙?�����Y�U���׶��..P0�("���:�^�eY� �d/J8��G�Yn�W"OOO7����?�m~�#y&���e`-Yl��"�e�J�@0%ˆ륖
^}�y�W��L������������3���������\���ja��-�V����p#I�T�t��'���G���~�W������8��e��K�O!��}2Q$��y
ټC�f��Qv-QhAmm_WϹ ~����l���xB���PY�U�����!_-K�M���O��b_��P���.b���C�\�zJ��{<Q�4,��×*�j�rwr��lk5I���l�&���hn^�T!� E�%kh �?`;�9���1H��*'(L,-#&�u�.%��)婒eB����^�5;�b=������:f��++�h6u���bq��u��q�x]�����s�wGw^����{�lC����T��Gqa:>o�~I [���[���p�6���%4�+$���=va���:s���!���"!h��m,�@�8�'?���N��z\��b�m�#O�O��;#�D�� �%� ^a�`"X�z�Ћx삳����7O�����:�B���_c;ÔQ���k��٬b{w�%����NCj����g�Xi��>����a�;�̡!qh���^���'w� �C>s��h�Y���`Y�ܳ��eE����))�x�ϐ��t��Ƭ�]��a�.�B��ߍoX��;I#����������&Iҡ��қ�.�։��j�*���S�g�Vo�Aw��Cx�Dx��Q�=�ŒZ��9�z�O���}�f����ܩ�tu*�x(ԎY	2�����!�"�pa,1�39:��
�v��͍��D!�B�������$��Ѝ����ښ�
�Eb��d������$Yф%1����@	��:]a�u���5��Yiv���3�6E$/�b��/3#�kK(o'+�)[�Y�#s�1qu�/r�D���]���dFw�s�m��Eۮ�(�(
�gͥ[����c�u����nF�bҐ��F̥�Ʒe�o2��"Z"�e�.�58�֛�LN ���њ9{�o�"?Sҥ�9ت*����åk��$���s㡤k�n��5�h�~`�4�E�'��΂�N\�C�7}��e۰2�j;/d�Mu��[��ѩ����C��a��l&<�o�nq8�Q��R��rm�x:{4T�8�.�w�u·,>#������O�sg��|�|��6{S�z���W!�̨��QH[�N��ZЮY��9%�/�}c��N��\��eL	q��ڤ��sL��/F%7&�9�#U����s�0�Kp���<��~��c}�7߻J{z�ș�0&��>�пg���P�M%o	\��_�a)�Q^Z�[�xt��`��9�+���y�j冟~FW��T��������Č^g�Yx �`OV�BVT����|� �Qc1�j�2E.G�ڽ�D�ݑ�eW+C=�u`�7OlYJ���m�\"y� �\�qOOZ�Zy4���X�V���q.��������&'J��bݥ�˝�r�$�H��a���W�h�q����}�5Ѫ;5��D`v�-�(�9S�,ҋD����8md���94a:cL5k�v#hr���	�lY�(z����$�X��zJ�}kl�mY۱FgQrRxC'�i�j�}�k�7�#1}X�-k[���$����S?����8m�c�P쳖�/�rE�hE�z0�`Qΐe�T �jq��bbu����S�pn1�y��es����ï���,��6��l�4�u�±޹<���k�	�<�"��(�8������7s ������(���,�B:�Z�V��8��ā;��/
g]�\�	�=�Z�nT���9ު��3��2E��XQ����
S]���ܨ�sP=���`�2�����Fw�!�h�6�Ro�su��4 +��cw�V��WWG��:Gc�ː�t ���˛��	���?2�n��k�ٶy$�g.����^B�F�T,�I ���6�����+Q ��G��(���odn%�Ⱥw;&�c�S�����˥�!�wq߲�t@V2���-�9�h�3���3��`nY�g�wy����m��$]��wN��X�b�_���/�-1p5�#3�8��mw�PӒ?%ٿڍ�!V$�,)��iAͩ�FW���X��	��g���r�(�"1�tvO�4�N�sH��Z�2&�bY�Ml�\p��8�A�w�>�o� *�I�"�8�_M�#������&<�����>S&�4��'������ݹ\^dbno%�!h����� 7�#]�W�L��a��P�pH��0��\�d�m[_'���Z����i�ZH�[91""�O��B' ��gA��O�=���Z�/�L�t�q�xH�������E+��j[%:��gn=�(�Z�T�Um*��:z�p��8�cpH�m�ĀY���/ұq!|]�n�T�u:c�~�(�4��1I��{�o�b"f^=�lEbH�U�7�����"�nk� �tj,P�W�x�+�������D�(U�
i���9x�q_&=&�U���j��+�p��ɅM�i��!��LW�Ѡ�N��])���f�e�@�7�І!Idp_�L'
���1�W^o��Yy��e�m���?��>j����ESR�$����Exu�,�pf���^X321]-�t'0�|��!�q̝W��9o#X���g��w�NNƖ�S�s�s����_��E��4�+�� � F��8YU�ZSS�b��Udʟ�!p'�	��B���jtk�liפ�3Y�a)��Q�ȑ���)���l�P�e#�s|1ݥv�|(���pd˭��C�ף4e)c�����jz�������ݽ��{	���2[?	����)rw��ާ ��q�%�.�ŞcCگ��R�z5�Uj��#S�u��΁Uj�MZ�#R�������\�ǡ)OO�!@G�eu^6����P>.�"��
-����R^��_��* ��h�v&��N�3�r���ڍ����{�C��^�<�k���p���2ؕ��~D4I{J�� )��aL�V�}'G���#���O�05��6����c���Q�ϙx{g�U��ࠚ[Z�� D�K�I\-Z�_�Ga���
)��"8��.\w�{"5���!R��_�6����ҭw=�N:�'=8�F���}�����\����'������	������s��D�P�SR*XQ"K�;����.�+�y�T������E�UO}����[�����[�[�O�?�
�M���d�R� T	y�+�8�j6�-�^��j�CT�H(7�������Po\��f>��[of�GBL��Mră7�.��sR�u=Wi���	�K'�Q���C�%��Yh�����,��w('���~���r���EɧO����(32�V�
]o�J6��{� ��Um�����?f���]���nұ!vTSB���P�^���s\�����}�p�"�>ܾ���m����@�g��>��P_����=V�'w�M���7���lK�X�ؙ��J?�f5��.�m�2n`�͐r���89���DK�պN�ء����~{�BOe���k���u�9d��cn��%�㖍g[�9��49�ȿKK񃻻�QQQ廤�=5~�C}��Y!Rr�h���3V�[��͎k���${^݀�Rp����([52Q�j���?T-X[��w�,�"��=���dEZ\\���0��K�i1�����I���>�Wۢ����0U�D�j3!�3�>e�l<�B%W�v�~	�D\>��ַ��Z�JϪk�@Ғ[G�i{��⒝���ԖG�Z����W��(7QK‾q�
�ȡW�.=k����QN��ƞ�Ƿ2��g&1�w�ѯX� ��:O�w
���	qފ
x�l�
Ƞz���^d�;�U��r��R�{���Ln���};����tz�j��wf3=w9}� [:;'655eEc��gffBD"�@���8�(�Ѹ\64�UЋ��ަn��u��_8_4觋�=�;�C� $HL+&P�{�KJ������6�,t���}%�#a#��\��i��@�G�����U�5��V�;���'�/��1�F��O���0~�u�]�-@�!C��M�A��=7�AUĎ���&$���H�DH��%��EJu�'E���hm��� b��n��\g�r!��2B�6��b�J%�H�X%�X�Y/iUlE1I����(�qm�A�O�\�3�b4��nUpݔ�GzؖK����� b�2 z�i����^�i�$QJ�.A�R�*��Lc���qf�[�F�j�Q�TH�A�n�U�c�C����	���)�0��P`:u���t�v	i����b�R�E�Ӓf����}X�����4�X�*JlW�.�0-��d�_d}}����#�x�	}�Qj��-g��%��o�[���C����2t��^-ځ�ǃ�-��D��4M\�ʄ	�]�ڨPkT�T���Iӈ��1�� {_��:��"M�:��R������v��=3�b4��	���rU�@��#��h��y��@;Ƕm�l��q1	T*ayyY�.ʀ��OS\ۄ�v���'
#�E�eI�0���׫���T*Ah��s�q0��!���:����B}�h�PVȃ�����l�a`����^����ԛ�\�pnFQ?����o��?����q��M;sĉ$#l�D�*ި�.j5����dr���o|���2á��Yaw�F�R�Zj`U��kgwHeH�^%
�*��j���ʏR^� ����T*�!X*[�u���������n �R)���O���[���`yyY	(���.+++DQDw�W�7)%�dk�:�e�x'1�SƮ9XV��q��0���E�\�U�LS����U$�{��#�u��Ϲ諸U�o��G�D�E�E���3�ʱ�1��$���$�^ل&�&�"@6Y8�d0�ăh�I&�c�2,�{L�"m��~UU��>O�ۗ4�T]�
� |4ϭ��s����}F֓�#Z->�+��e�֤���zY��EI��k�Z�^��0�p]�;w�G?�	��/}�K�~�"wn�&�)�i�c�ʏ�7=B�R�0(�H�L#k�?B&�c	���7�Z	��m֏��?�c,L��0A�HbI��yP�F��D�S��K鯞8A�QG�U�ya�4}�q.��aN�(��u�I�w�!�t����ȉ�8�J�G���p���40=H5A���[�6#)�	�j�1�ZI���z]ͤ2��޻Gݟ��H�n"�4U�2ɖnt/F)RJD����f*���x<ƭV�Tk���U.5�ط�!��O��.}�W?����q��]�F*��G`�T*�Iİ��^�id��\?WG!�n��O�������'>�������m���$XB>�U��	`96q�0�#66_�0>��#����kTj5Z��X�	P��.&�_������&.\��T�	'gΜ����� �kд1�uj����]\���5^z�%�߿��%�vU���l6����������ɣ�>*���0�a�!V���;C)C��+�A
��x����/�������	���p���u��Y�k �m�L%�h�1��0O���((�I�`}�{�GKV��y�3�4��#N�<�L-�j5���}~%���eBO�-􆋬�B@G����r��I����nﳶ����"��V^w�m[	Ogan11W���J�QC��2T����&v�S]~�g/�η��J�?%'��B2hu	{�c��wh��sok���e�c�� ���6�qH���N�����9���Z��NP�I3
���F˶��gϞe4�7�8?u�~]MRk�����P��y��wI��Sm#!��1
�DA��)�s'wn�18�2F׭�oY,/���ɂ����AL
� L�D���2Q�k?f��o1d��8��WU����*�7_ckg�ᨏ_�9~�87o��kIE�0}b��a��eZD���BR$/��"պ�aܼy��/�b�)�x�iC旚[��؂PJ���?��?�Fw�E}q1��JS���}��a� �a<�a�ק<<%�[���1���M���>�0J�Z��ܺu��}���0vk	�2��lp��\�r�o����B��;ɘ4M�Pi�����2���S�c�;V�IV�W�� R*��f�cǎ����o����eww����4�ƃ���vH#�(ngo�V�E��֔��:=V��4M� ȣ;=���\�É9!�c#b���_�9�u�V��a����2��I�6�iX�Q̉��p �6���t��F��82�	v���ؘ�E�WM�K�����gz��Q���̻ex!)�L0=��8h��dt�8Qw%��!z5�{w�x�w�8w��u�kN�P����y�p�{׮���!��2�0D&	�e���`��J1
9���� �˰iz>{w��̨�	�шz}� �#N?����.B*
�h4�G���cG�qC�a��!v�F�v��k��`���O���2Mj5���}<����$�%/.����-�����V�E�9�p<���3�;-^|���9�����C��0BP�}���XXX��HI!�j[T���R�$������Ǹw��/���w9~�,����I���p��9��ܾs��AhJ�~ �6��v�� ���H1<�B	��TeA
HD69]�}�fD� �b,�����W���A�94��*X��Ƶd�V�0��Fܹs��8�>��I��4�sz�Ƈ�oߧV���UfZ�R�!�l���Kc��G7>���$���l�ߺO(G���,L��a�)�r�������GW����]���uKU�ۭ��q�zD��iS��Y=��ضK�a2��K������������v�o��t9��
g_}����g+�z=�D��秋��&RT=�,�$�0T�F�������4���9d0���+�� &��D��	�_���[,--������I��n��1 ��K��,��F�US�!�>�i����:[�c���K���a���UH�'��,�y�j��e�� ���_�3�}H��� �0�"bէ+@�b`H�Ȕ�D!�4b�s���2?��x&���&�%	��1̔4U����/h�]n߹A��2�p�����$2&��B�����1�G�������.�N�I��ģ�������txU�URo���wh��BQ=�]����4���w�JBFq����I�ʢ�:�,�J�cm�8?��2Y�ۘ{�昛���'q�):`�)],�Cn��(���XY�N��ad�Wf���Tƪ�t��F�.����m3GHT�EA0���f����z������j��=��m`��,4�$��4I��$���H�È$N1��t8y�,���"���[�ܡ}0��X^�(6�1�tq�
�b���G]�$ �F��T��>�h4bgo)^9�*����%��N�K%$�Ķ�<l�!�$!����7	�1�q�51��Li�����dnn�n����6RʼH�����y9(�1a4D	�a�Ѩ�0b���[��s�c�YB�D�iILK�7n��f���-��:��~���$ID�D�1$���k�쑪�I�5���|R��xj�
X��EE=T���j�
�_�%<� RSҬU�l�A�mJ\��6!�c��׳�*��K��v��yY.����Q`�:s|�w�k�^f��݃��P`ul�Ǳ�Xf��iT�z��5�2����D%�eR�UU�!�ٕ�벾���ٗY\^�Дǜ�!����\u��J�e4��u{�j5�{�.��ַ�F�͸B ����8�1�(P�L�ƶܼ`x��/�T]N��b�)q2fo�>�/�´���R�T��eY�|�q�`����p�K?���:T�l��2��EF7�lLS��	Q��:MS�ՠ(#Q�K�$���01-A'��,�[3����<**��:�T󾑒�RI�][t����矪� �ǲ��Yẖ�����0"�b�PҘ[B
��p��۩0����`��L�ڜ���a����q�iݧ�8�A8HeB��!�z}u�۶M��Y�'���n�ĊG3X]=�������ͫխV������9??�A��@ɣ�贈a�:��`6F�7�礔�Z-�x�HF��׿2��pH�����ܼy�S��8P|�̉ͯ�ܕ�ٵ�<�����5��2U�XH�8�ÀJ�J���v,�z��(�NZv�T-<�i
Q4"�TVP�{�4lR�湕�|i��B���Klݾ����9�c�峸F��[}l���m�!�2?�Z������>O�V'�$����%G���s�4�sj�H1����{�߻����4j>�c2�P��g��kS��H���TB�|N���1++6+++�޿��8��ѣGsy�;w��.+++�;w�q�
U�6ۖK�L,K2���-s�����t:��y� �s�������n��ƧO]��u�~oĹ��z�a�H��:nN��l[}�˗/�^W�{}nݺ����HŘ�*V��ނ8���k9yZ��:�f�X3��X���F���͛ԫ1/\��n������S~����&�pY\XQ�f���쯔�P���z$���>���5VWW9v�����4}��6�v;�^����
���[ �Y�e�Z�R�Jƣ�h(f���D��&Q����N���S�n�z��F�dIν�]�����v�
A(���x������aܦ��c�����>��D��~�j�Ā�Ԛ��~������f4R�`0ȧ�i#y؀�X��:�Mm�L,JPmԱ��u�$I�����3�>��~�ߔ�����,/]�$/_�,/^�(�(�:��>�}�������[��ߺ,��w�ȗ_{]�˷ORNl�k׾��s��/|��W����߻��z����oO�3=.� �j������<	^{�?j4���������;�v��Y}��B�[�7����"��Z��'������t9�14EG��U�xAzk6ڤ��3��Y�O��6��!�Φ��bW����IF=.tw@�Z��ޫg�O7n�CWpA�0��hFГB���*	�XtΦ�N�1��Cu��8.�`4�L�rt����?K���9-�i�)� ��/Ӈ�\�"?��ʳ��u�u�i��<�@��|�~|Ys�'��5����܇�vv��L�T�6I<y�X�h4Ĕ)�2cF!�����c��2�L�p�ö��5Mϓ<���3�?I7ߓB��گ�$݅O}�i��+iB�WB���F�C����_��ѓF�����ӂ�y�'���:oQ���Mjp��U���d�b��`�w���+���(s=����"s�(vk�y�>.f�`,��F����5-B��M�T4�	C���tiL�=t]G'�tޢ,xރ�f��`�t�g13-�i��Ρξ�Y�z��2PJfY3�����,0����nPj��0m&�noH�H�p�d%�dE	�Wͅ��3m0:��=�A���:�C��&Cj�Z.SV�:�h]�g��vzu�5�_Z�h-��0J���Plڟ��	�qNd�|�2�� ���J�d0��<&��.���3m0Z�R��U=ֈ�z���U�?�ӧOO|�(��̴��n<}E��Sh�kOw ���o��Ǆ�uc�4�03���nY6f��W���M]�Ų,�޽K0����z�k��;-����Lk�l�n���{/��8I��\qt�N�q��Fy߰���}�����!�b�0±l<�x�^�4A0������Z�D��uϗO�.�tv���t���u<K��	S��)e����_�%e�Q�r�3m0�J�P��8U�$�om4zz�$�O��h��`&�z�^�����VY�i���1ד�'M��G�>z��iF��$�j]u]���ݯ�փ\�xTO�i��a��O<7�	A-+�/h�j�}�a�M�,�+�̴�茫�*�C�ȅ�ҒjZ�p1�>���6�l���~��َI�q\�$I҈2*I��*91%O6-��'yB���Q�y�s��he\��|ӆ�7��Tٲ�z���T�CZ,uLf�`tۇ*z�vQ��LL�3�Sa\��|x�DYT�� �i�LGI �j� �0�J/h�E'��q����J~��	�Cв����E�0�8cjҘ��G��?a��>�a����wp���ӥ��Q�!�3}�h����=�Q�$���B�R��Wq]�4��a�ӂ�6-������u�Hk=��6~Mݘ�|�L(�W;�e7�۶��6�b�g�x8���`&�^����j��Xf�,�7��O��&��Sa�(�L[�z�f<s���|tr��I�tY�ƓEc�Ʋ�\��i�B�ϭ�8e��E����3m0��q�����=_d��碈��է���h�vL�x�������L'���T�yQ�l8����H5����N|}���OZ�L��>j��m�Ξ�SD,˿(J�=�a&�ZM���ɢ�#�25t�u�i����I� �^����2�h��8��L�4(t>7�	a8�Uc����� yBM����Q<jd��L��ԽBOÇ�b�_���)NK�&c�78=u{i��#���&���OSY f�`t-GJ���j���H����2	�3m0�b�ia�-֏�c%�����ۍ�m�p��ɈJ�"�4������������Y����+˼x�%���Q�k�A�Z����f���n{�k���s��ܱ�<�k�{��<	f������5N��N�&��8^�z���_=}�4������������f)kmllP��B��/|�Ry̜�H)���R޾}[�axOX&�mq��}�%ʕ���u��666�p��i��o"��:�u�A.�����7���JS�x\�ԕ4�|�0�Vw���2��VJY.BGb[[[�qL��accୌ#3����H����}��$�ˉafN)�Y���E��u����V��S��8{��gΐ�db�]JyU�2Ǖ+W���G���\�t��p���oI)e�2�cY�'~)��R&��������ŋ'�q>5��W�نJ��y    IEND�B`�PK   ��U�0�	  �5     jsons/user_defined.json�Zm���+}^g����F۠I��i��0
��l�骓j��{�|wN��$.�/��!�|ކ�O��ǻ~�br��w�Z����_N�����z��/����ü|�~�⟟������ݟv��j���~�����]������#>;�+
߼�R�m7Y/���yO�4���H�0�K�Ӡ�Z�_̣ϨS&����ݡ�ƫ�~�[����<�?��ww�w���z��f����4�~~�����}|���sN�)�>������WA�x���â6��0��w�7���z���u���[��bvB�.9O>
>���f�x���ۏOz;������zy��l���������oo�NC��C�~����#�`9�F�;�&��7�@X�7��m���~}�n�b��&e濆����p��w���0��S��R���~55Z�e/=Q�# I� �����xs!���/�z�D�o!�6��t�_����%�bg��/�@�s��S��?�x����a��nn~�.��%`\��rI3�>�r�V��ij�ł8��<�G�����<v3q��� ��ԀF��BNA:I s<��7�w���5�<?�(@&��~ /��! �{}�_�k��kP�����VӴ����ibIS]e�S�W�y*/(	*�S�UT�SJ$�@|p�$��]����5,_���+@�� )�`*�@/���n���,g��a����a��y�^��o?N��7��g�����x��?����7�gK��K����~)��m� ˜�im
��I�h���^R�{��-�	Ee
�AQc 'f>v�Q��ᷱ{nc2G9��x��Ѳ?�k�=&�O����z=��W�XEr���]6�Z=�C' Au)�H&m�.���pؤF�nx�ɷVס���2�Oi@�"7����3vU� Jɚ��A�,� %sG��@E�\sr�zʨ����a�&%�;��ȅ@�C&Gdg����C�2"r�>iW�ęGRh.?�k�����%�Jع��z��,���`m<lA?�O~H�c.�$�-����ه��++�����Kn�}��ǥ��!��X���Ǌ�@ ���DR��f\Ɗ����N\ʛ��Ξ(�.?Th�3A�	�*n,�+}Er��b� LV�
��,Ʊ�9���-6II���T­O�X�����M$7ׯd[*���A���
�S��+�6 ��M~0C3nW5�o)��a�9ñ���K�!i���9y.���?��HT��]J�!�R��u�-4��+u9��a3����H�x��Aq0������L�A���H;�!�r4�A*����07��*���;��eh�7'�����+����XV��+�1Rw4�eC&�Ծ�^QB�͑Jځ�iF�y��� U\k�.��� �t�DBj�O�������`�I$��n��e�$�!����m����X� ]�������BT����E�������^}�[9hk�&pC�Ќ�Tc-?��X�dҞ�+=D�]��K���q�*]x[�McԢk�>0j�j����c Q���}���'΀Nʀ`��%#��"=��a*�}"ӈ^�*��Y���%*M#l�=�Ňbd�n��*�ə�ӡ����%�Kj p͡�T9Q����Vb�:�C�}&����0�NS H=7�3UR���	����%�� �hL�B����/�#��`��* ��B(qj$.%��%M�%J;B����,CF�o�g�Q�l��Cv�����kOmo1ݘ�1����ĳ<��q�΀��h�T���"��6Dɸ$8R�%1@��Z0j�� a��r�1�Mљ*�M��h�d|�r�'�	Z�D�=��,�?1��;������W�IO'z�.$�v}����xN:�}��l�}�\���>w�޴d�fn�ğ!�C�i�^M���|W:�L{gW�~H����Ͼ}kk�/X��Ύt>�yk�_����?^�|�V�$��a���15kNM��:�m����@�vѬ�~yw�xlR^��Ͽ&����5����4q3sk�tj��F�4��/Ek̅����0��Bܼ�\an9�F��ԉ������\�`CW�\ry�\��\d*��FN"�3���M�Z4?�_B͆�5�UdCn;j��sr���U<Lߠ��lr�jr����;il��&�!?q��f�Xa-:�8��Q�Gu���Z��p�J����k�N�Ѷ�`J�E������z�c�f�c�K��o�*�/��s2�`;h'�%Sj��e��X0,Z8{��t�Z���j>��jZkR�8X Byմڢ�"�LP�'UZ��ǣ�r�ɍ�i�ܛ=�#�*p;�bW��~���C�Ɉ�W�
������WjWd��6s.���Q��J�[�*k�B�f_R8�k�k��k�S�M��v/Oõ>!*@s�"����~�?\|��k})���wq��b�Su=ug���OW�����7/^�k�^|����Ͽ PK
   ��U܌W�Sq  �                  cirkitFile.jsonPK
   �R�Ts�7+5J  dK  /             �q  images/6c71542d-16cb-4630-930f-71c4de5e1144.pngPK
   �R�T��4�� ̻ /             �  images/7a4be1c8-201b-41f2-b584-263fc50cb409.pngPK
   Y�U���@Y�	 �
 /             8x images/8464ed5e-37c3-43b3-8b47-7240858568a5.pngPK
   �R�T��K� 	� /             �T images/cd1eebff-8d4c-4172-8358-6f93b12ef793.pngPK
   �R�T��!�D�  Ԟ  /             v� images/cf2dd1a8-295d-437f-92b8-7fcc138ae9be.pngPK
   ��U�0�	  �5               � jsons/user_defined.jsonPK      S  �   